// nios_simple.v

// Generated using ACDS version 13.0sp1 232 at 2024.03.29.14:49:18

`timescale 1 ps / 1 ps
module nios_simple (
		inout  wire [7:0]  tri_state_bridge_flash_data,              //       tri_state_bridge_flash_bridge_0_out.tri_state_bridge_flash_data
		output wire [0:0]  write_n_to_the_cfi_flash,                 //                                          .write_n_to_the_cfi_flash
		output wire [0:0]  select_n_to_the_cfi_flash,                //                                          .select_n_to_the_cfi_flash
		output wire [0:0]  read_n_to_the_cfi_flash,                  //                                          .read_n_to_the_cfi_flash
		output wire [22:0] tri_state_bridge_flash_address,           //                                          .tri_state_bridge_flash_address
		input  wire        reset_n,                                  //                      clk_ext_clk_in_reset.reset_n
		input  wire        clk_ext,                                  //                            clk_ext_clk_in.clk
		output wire        pll_c0_out,                               //                                    pll_c0.clk
		output wire        pll_c1_out,                               //                                c1_out_clk.clk
		output wire        pll_c2_out,                               //                                c2_out_clk.clk
		output wire        pll_c3_out,                               //                                c3_out_clk.clk
		output wire        locked_from_the_pll,                      //                        pll_locked_conduit.export
		output wire        phasedone_from_the_pll,                   //                     pll_phasedone_conduit.export
		output wire [12:0] zs_addr_from_the_sdram,                   //                                sdram_wire.addr
		output wire [1:0]  zs_ba_from_the_sdram,                     //                                          .ba
		output wire        zs_cas_n_from_the_sdram,                  //                                          .cas_n
		output wire        zs_cke_from_the_sdram,                    //                                          .cke
		output wire        zs_cs_n_from_the_sdram,                   //                                          .cs_n
		inout  wire [31:0] zs_dq_to_and_from_the_sdram,              //                                          .dq
		output wire [3:0]  zs_dqm_from_the_sdram,                    //                                          .dqm
		output wire        zs_ras_n_from_the_sdram,                  //                                          .ras_n
		output wire        zs_we_n_from_the_sdram,                   //                                          .we_n
		output wire [23:0] RGB_OUT_from_the_video_sync_generator,    //                 video_sync_generator_sync.RGB_OUT
		output wire        HD_from_the_video_sync_generator,         //                                          .HD
		output wire        VD_from_the_video_sync_generator,         //                                          .VD
		output wire        DEN_from_the_video_sync_generator,        //                                          .DEN
		output wire        spi_data_out_from_the_sd_card_controller, //    sd_card_controller_avalon_slave_export.data_out
		input  wire        spi_data_in_to_the_sd_card_controller,    //                                          .data_in
		output wire        spi_cs_n_from_the_sd_card_controller,     //                                          .cs_n
		output wire        spi_clk_from_the_sd_card_controller,      //                                          .clk
		output wire        out_port_from_the_lcd_i2c_scl,            //           lcd_i2c_scl_external_connection.export
		output wire        out_port_from_the_lcd_i2c_en,             //            lcd_i2c_en_external_connection.export
		inout  wire        bidir_port_to_and_from_the_lcd_i2c_sda,   //           lcd_i2c_sda_external_connection.export
		input  wire        MISO_to_the_touch_panel_spi,              //                  touch_panel_spi_external.MISO
		output wire        MOSI_from_the_touch_panel_spi,            //                                          .MOSI
		output wire        SCLK_from_the_touch_panel_spi,            //                                          .SCLK
		output wire        SS_n_from_the_touch_panel_spi,            //                                          .SS_n
		input  wire        in_port_to_the_touch_panel_pen_irq_n,     // touch_panel_pen_irq_n_external_connection.export
		input  wire        in_port_to_the_touch_panel_busy,          //      touch_panel_busy_external_connection.export
		inout  wire [15:0] SRAM_DQ_to_and_from_the_sram,             //                          sram_conduit_end.DQ
		output wire [19:0] SRAM_ADDR_from_the_sram,                  //                                          .ADDR
		output wire        SRAM_UB_n_from_the_sram,                  //                                          .UB_n
		output wire        SRAM_LB_n_from_the_sram,                  //                                          .LB_n
		output wire        SRAM_WE_n_from_the_sram,                  //                                          .WE_n
		output wire        SRAM_CE_n_from_the_sram,                  //                                          .CE_n
		output wire        SRAM_OE_n_from_the_sram                   //                                          .OE_n
	);

	wire          sgdma_pixel_out_endofpacket;                                                                           // sgdma_pixel:out_endofpacket -> timing_adapter:in_endofpacket
	wire          sgdma_pixel_out_valid;                                                                                 // sgdma_pixel:out_valid -> timing_adapter:in_valid
	wire          sgdma_pixel_out_startofpacket;                                                                         // sgdma_pixel:out_startofpacket -> timing_adapter:in_startofpacket
	wire    [1:0] sgdma_pixel_out_empty;                                                                                 // sgdma_pixel:out_empty -> timing_adapter:in_empty
	wire   [31:0] sgdma_pixel_out_data;                                                                                  // sgdma_pixel:out_data -> timing_adapter:in_data
	wire          sgdma_pixel_out_ready;                                                                                 // timing_adapter:in_ready -> sgdma_pixel:out_ready
	wire          timing_adapter_out_endofpacket;                                                                        // timing_adapter:out_endofpacket -> fifo:avalonst_sink_endofpacket
	wire          timing_adapter_out_valid;                                                                              // timing_adapter:out_valid -> fifo:avalonst_sink_valid
	wire          timing_adapter_out_startofpacket;                                                                      // timing_adapter:out_startofpacket -> fifo:avalonst_sink_startofpacket
	wire    [1:0] timing_adapter_out_empty;                                                                              // timing_adapter:out_empty -> fifo:avalonst_sink_empty
	wire   [31:0] timing_adapter_out_data;                                                                               // timing_adapter:out_data -> fifo:avalonst_sink_data
	wire          timing_adapter_out_ready;                                                                              // fifo:avalonst_sink_ready -> timing_adapter:out_ready
	wire          pixel_converter_out_endofpacket;                                                                       // pixel_converter:eop_out -> video_sync_generator:eop
	wire          pixel_converter_out_valid;                                                                             // pixel_converter:valid_out -> video_sync_generator:valid
	wire          pixel_converter_out_startofpacket;                                                                     // pixel_converter:sop_out -> video_sync_generator:sop
	wire          pixel_converter_out_empty;                                                                             // pixel_converter:empty_out -> video_sync_generator:empty
	wire   [23:0] pixel_converter_out_data;                                                                              // pixel_converter:data_out -> video_sync_generator:data
	wire          pixel_converter_out_ready;                                                                             // video_sync_generator:ready -> pixel_converter:ready_in
	wire          fifo_out_endofpacket;                                                                                  // fifo:avalonst_source_endofpacket -> fifo_to_pixel_converter:in_endofpacket
	wire          fifo_out_valid;                                                                                        // fifo:avalonst_source_valid -> fifo_to_pixel_converter:in_valid
	wire          fifo_out_startofpacket;                                                                                // fifo:avalonst_source_startofpacket -> fifo_to_pixel_converter:in_startofpacket
	wire    [1:0] fifo_out_empty;                                                                                        // fifo:avalonst_source_empty -> fifo_to_pixel_converter:in_empty
	wire   [31:0] fifo_out_data;                                                                                         // fifo:avalonst_source_data -> fifo_to_pixel_converter:in_data
	wire          fifo_out_ready;                                                                                        // fifo_to_pixel_converter:in_ready -> fifo:avalonst_source_ready
	wire          fifo_to_pixel_converter_out_endofpacket;                                                               // fifo_to_pixel_converter:out_endofpacket -> pixel_converter:eop_in
	wire          fifo_to_pixel_converter_out_valid;                                                                     // fifo_to_pixel_converter:out_valid -> pixel_converter:valid_in
	wire          fifo_to_pixel_converter_out_startofpacket;                                                             // fifo_to_pixel_converter:out_startofpacket -> pixel_converter:sop_in
	wire    [1:0] fifo_to_pixel_converter_out_empty;                                                                     // fifo_to_pixel_converter:out_empty -> pixel_converter:empty_in
	wire   [31:0] fifo_to_pixel_converter_out_data;                                                                      // fifo_to_pixel_converter:out_data -> pixel_converter:data_in
	wire          fifo_to_pixel_converter_out_ready;                                                                     // pixel_converter:ready_out -> fifo_to_pixel_converter:out_ready
	wire   [22:0] tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_address_out;                             // tri_state_bridge_flash_pinSharer_0:tri_state_bridge_flash_address -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_address
	wire    [7:0] tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_in;                                 // tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_in -> tri_state_bridge_flash_pinSharer_0:tri_state_bridge_flash_data_in
	wire    [7:0] tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_out;                                // tri_state_bridge_flash_pinSharer_0:tri_state_bridge_flash_data -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data
	wire          tri_state_bridge_flash_pinsharer_0_tcm_grant;                                                          // tri_state_bridge_flash_bridge_0:grant -> tri_state_bridge_flash_pinSharer_0:grant
	wire    [0:0] tri_state_bridge_flash_pinsharer_0_tcm_select_n_to_the_cfi_flash_out;                                  // tri_state_bridge_flash_pinSharer_0:select_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_select_n_to_the_cfi_flash
	wire          tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_outen;                              // tri_state_bridge_flash_pinSharer_0:tri_state_bridge_flash_data_outen -> tri_state_bridge_flash_bridge_0:tcs_tri_state_bridge_flash_data_outen
	wire          tri_state_bridge_flash_pinsharer_0_tcm_request;                                                        // tri_state_bridge_flash_pinSharer_0:request -> tri_state_bridge_flash_bridge_0:request
	wire    [0:0] tri_state_bridge_flash_pinsharer_0_tcm_write_n_to_the_cfi_flash_out;                                   // tri_state_bridge_flash_pinSharer_0:write_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_write_n_to_the_cfi_flash
	wire    [0:0] tri_state_bridge_flash_pinsharer_0_tcm_read_n_to_the_cfi_flash_out;                                    // tri_state_bridge_flash_pinSharer_0:read_n_to_the_cfi_flash -> tri_state_bridge_flash_bridge_0:tcs_read_n_to_the_cfi_flash
	wire          cfi_flash_tcm_chipselect_n_out;                                                                        // cfi_flash:tcm_chipselect_n_out -> tri_state_bridge_flash_pinSharer_0:tcs0_chipselect_n_out
	wire          cfi_flash_tcm_grant;                                                                                   // tri_state_bridge_flash_pinSharer_0:tcs0_grant -> cfi_flash:tcm_grant
	wire          cfi_flash_tcm_data_outen;                                                                              // cfi_flash:tcm_data_outen -> tri_state_bridge_flash_pinSharer_0:tcs0_data_outen
	wire          cfi_flash_tcm_request;                                                                                 // cfi_flash:tcm_request -> tri_state_bridge_flash_pinSharer_0:tcs0_request
	wire    [7:0] cfi_flash_tcm_data_out;                                                                                // cfi_flash:tcm_data_out -> tri_state_bridge_flash_pinSharer_0:tcs0_data_out
	wire          cfi_flash_tcm_write_n_out;                                                                             // cfi_flash:tcm_write_n_out -> tri_state_bridge_flash_pinSharer_0:tcs0_write_n_out
	wire   [22:0] cfi_flash_tcm_address_out;                                                                             // cfi_flash:tcm_address_out -> tri_state_bridge_flash_pinSharer_0:tcs0_address_out
	wire    [7:0] cfi_flash_tcm_data_in;                                                                                 // tri_state_bridge_flash_pinSharer_0:tcs0_data_in -> cfi_flash:tcm_data_in
	wire          cfi_flash_tcm_read_n_out;                                                                              // cfi_flash:tcm_read_n_out -> tri_state_bridge_flash_pinSharer_0:tcs0_read_n_out
	wire          cpu_instruction_master_waitrequest;                                                                    // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [27:0] cpu_instruction_master_address;                                                                        // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                           // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                       // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                                  // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire          cpu_data_master_waitrequest;                                                                           // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                             // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [27:0] cpu_data_master_address;                                                                               // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                 // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                  // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                              // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                           // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire          cpu_data_master_readdatavalid;                                                                         // cpu_data_master_translator:av_readdatavalid -> cpu:d_readdatavalid
	wire    [3:0] cpu_data_master_byteenable;                                                                            // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          sgdma_pixel_descriptor_write_waitrequest;                                                              // sgdma_pixel_descriptor_write_translator:av_waitrequest -> sgdma_pixel:descriptor_write_waitrequest
	wire   [31:0] sgdma_pixel_descriptor_write_writedata;                                                                // sgdma_pixel:descriptor_write_writedata -> sgdma_pixel_descriptor_write_translator:av_writedata
	wire   [31:0] sgdma_pixel_descriptor_write_address;                                                                  // sgdma_pixel:descriptor_write_address -> sgdma_pixel_descriptor_write_translator:av_address
	wire          sgdma_pixel_descriptor_write_write;                                                                    // sgdma_pixel:descriptor_write_write -> sgdma_pixel_descriptor_write_translator:av_write
	wire          sgdma_pixel_descriptor_read_waitrequest;                                                               // sgdma_pixel_descriptor_read_translator:av_waitrequest -> sgdma_pixel:descriptor_read_waitrequest
	wire   [31:0] sgdma_pixel_descriptor_read_address;                                                                   // sgdma_pixel:descriptor_read_address -> sgdma_pixel_descriptor_read_translator:av_address
	wire          sgdma_pixel_descriptor_read_read;                                                                      // sgdma_pixel:descriptor_read_read -> sgdma_pixel_descriptor_read_translator:av_read
	wire   [31:0] sgdma_pixel_descriptor_read_readdata;                                                                  // sgdma_pixel_descriptor_read_translator:av_readdata -> sgdma_pixel:descriptor_read_readdata
	wire          sgdma_pixel_descriptor_read_readdatavalid;                                                             // sgdma_pixel_descriptor_read_translator:av_readdatavalid -> sgdma_pixel:descriptor_read_readdatavalid
	wire          sgdma_pixel_m_read_waitrequest;                                                                        // sgdma_pixel_m_read_translator:av_waitrequest -> sgdma_pixel:m_read_waitrequest
	wire   [31:0] sgdma_pixel_m_read_address;                                                                            // sgdma_pixel:m_read_address -> sgdma_pixel_m_read_translator:av_address
	wire          sgdma_pixel_m_read_read;                                                                               // sgdma_pixel:m_read_read -> sgdma_pixel_m_read_translator:av_read
	wire   [31:0] sgdma_pixel_m_read_readdata;                                                                           // sgdma_pixel_m_read_translator:av_readdata -> sgdma_pixel:m_read_readdata
	wire          sgdma_pixel_m_read_readdatavalid;                                                                      // sgdma_pixel_m_read_translator:av_readdatavalid -> sgdma_pixel:m_read_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                      // cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                        // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                          // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                            // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                             // cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                         // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                      // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                       // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire   [15:0] sram_avalon_slave_translator_avalon_anti_slave_0_writedata;                                            // sram_avalon_slave_translator:av_writedata -> sram:s_writedata
	wire   [19:0] sram_avalon_slave_translator_avalon_anti_slave_0_address;                                              // sram_avalon_slave_translator:av_address -> sram:s_address
	wire          sram_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                           // sram_avalon_slave_translator:av_chipselect -> sram:s_chipselect_n
	wire          sram_avalon_slave_translator_avalon_anti_slave_0_write;                                                // sram_avalon_slave_translator:av_write -> sram:s_write_n
	wire          sram_avalon_slave_translator_avalon_anti_slave_0_read;                                                 // sram_avalon_slave_translator:av_read -> sram:s_read_n
	wire   [15:0] sram_avalon_slave_translator_avalon_anti_slave_0_readdata;                                             // sram:s_readdata -> sram_avalon_slave_translator:av_readdata
	wire    [1:0] sram_avalon_slave_translator_avalon_anti_slave_0_byteenable;                                           // sram_avalon_slave_translator:av_byteenable -> sram:s_byteenable_n
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                   // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                     // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [24:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                       // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                    // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                         // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                          // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [31:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                      // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                                 // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [3:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                    // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_waitrequest;                                              // cfi_flash:uas_waitrequest -> cfi_flash_uas_translator:av_waitrequest
	wire    [0:0] cfi_flash_uas_translator_avalon_anti_slave_0_burstcount;                                               // cfi_flash_uas_translator:av_burstcount -> cfi_flash:uas_burstcount
	wire    [7:0] cfi_flash_uas_translator_avalon_anti_slave_0_writedata;                                                // cfi_flash_uas_translator:av_writedata -> cfi_flash:uas_writedata
	wire   [22:0] cfi_flash_uas_translator_avalon_anti_slave_0_address;                                                  // cfi_flash_uas_translator:av_address -> cfi_flash:uas_address
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_lock;                                                     // cfi_flash_uas_translator:av_lock -> cfi_flash:uas_lock
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_write;                                                    // cfi_flash_uas_translator:av_write -> cfi_flash:uas_write
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_read;                                                     // cfi_flash_uas_translator:av_read -> cfi_flash:uas_read
	wire    [7:0] cfi_flash_uas_translator_avalon_anti_slave_0_readdata;                                                 // cfi_flash:uas_readdata -> cfi_flash_uas_translator:av_readdata
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_debugaccess;                                              // cfi_flash_uas_translator:av_debugaccess -> cfi_flash:uas_debugaccess
	wire          cfi_flash_uas_translator_avalon_anti_slave_0_readdatavalid;                                            // cfi_flash:uas_readdatavalid -> cfi_flash_uas_translator:av_readdatavalid
	wire    [0:0] cfi_flash_uas_translator_avalon_anti_slave_0_byteenable;                                               // cfi_flash_uas_translator:av_byteenable -> cfi_flash:uas_byteenable
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_writedata;                                                // pll_pll_slave_translator:av_writedata -> pll:writedata
	wire    [1:0] pll_pll_slave_translator_avalon_anti_slave_0_address;                                                  // pll_pll_slave_translator:av_address -> pll:address
	wire          pll_pll_slave_translator_avalon_anti_slave_0_write;                                                    // pll_pll_slave_translator:av_write -> pll:write
	wire          pll_pll_slave_translator_avalon_anti_slave_0_read;                                                     // pll_pll_slave_translator:av_read -> pll:read
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_readdata;                                                 // pll:readdata -> pll_pll_slave_translator:av_readdata
	wire   [31:0] sgdma_pixel_csr_translator_avalon_anti_slave_0_writedata;                                              // sgdma_pixel_csr_translator:av_writedata -> sgdma_pixel:csr_writedata
	wire    [3:0] sgdma_pixel_csr_translator_avalon_anti_slave_0_address;                                                // sgdma_pixel_csr_translator:av_address -> sgdma_pixel:csr_address
	wire          sgdma_pixel_csr_translator_avalon_anti_slave_0_chipselect;                                             // sgdma_pixel_csr_translator:av_chipselect -> sgdma_pixel:csr_chipselect
	wire          sgdma_pixel_csr_translator_avalon_anti_slave_0_write;                                                  // sgdma_pixel_csr_translator:av_write -> sgdma_pixel:csr_write
	wire          sgdma_pixel_csr_translator_avalon_anti_slave_0_read;                                                   // sgdma_pixel_csr_translator:av_read -> sgdma_pixel:csr_read
	wire   [31:0] sgdma_pixel_csr_translator_avalon_anti_slave_0_readdata;                                               // sgdma_pixel:csr_readdata -> sgdma_pixel_csr_translator:av_readdata
	wire   [31:0] fifo_in_csr_translator_avalon_anti_slave_0_writedata;                                                  // fifo_in_csr_translator:av_writedata -> fifo:wrclk_control_slave_writedata
	wire    [2:0] fifo_in_csr_translator_avalon_anti_slave_0_address;                                                    // fifo_in_csr_translator:av_address -> fifo:wrclk_control_slave_address
	wire          fifo_in_csr_translator_avalon_anti_slave_0_write;                                                      // fifo_in_csr_translator:av_write -> fifo:wrclk_control_slave_write
	wire          fifo_in_csr_translator_avalon_anti_slave_0_read;                                                       // fifo_in_csr_translator:av_read -> fifo:wrclk_control_slave_read
	wire   [31:0] fifo_in_csr_translator_avalon_anti_slave_0_readdata;                                                   // fifo:wrclk_control_slave_readdata -> fifo_in_csr_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                  // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                    // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                 // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                      // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                       // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                   // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                            // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                           // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] descriptor_mem_s1_translator_avalon_anti_slave_0_writedata;                                            // descriptor_mem_s1_translator:av_writedata -> descriptor_mem:writedata
	wire   [13:0] descriptor_mem_s1_translator_avalon_anti_slave_0_address;                                              // descriptor_mem_s1_translator:av_address -> descriptor_mem:address
	wire          descriptor_mem_s1_translator_avalon_anti_slave_0_chipselect;                                           // descriptor_mem_s1_translator:av_chipselect -> descriptor_mem:chipselect
	wire          descriptor_mem_s1_translator_avalon_anti_slave_0_clken;                                                // descriptor_mem_s1_translator:av_clken -> descriptor_mem:clken
	wire          descriptor_mem_s1_translator_avalon_anti_slave_0_write;                                                // descriptor_mem_s1_translator:av_write -> descriptor_mem:write
	wire   [31:0] descriptor_mem_s1_translator_avalon_anti_slave_0_readdata;                                             // descriptor_mem:readdata -> descriptor_mem_s1_translator:av_readdata
	wire    [3:0] descriptor_mem_s1_translator_avalon_anti_slave_0_byteenable;                                           // descriptor_mem_s1_translator:av_byteenable -> descriptor_mem:byteenable
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                       // peripheral_bridge:s0_waitrequest -> peripheral_bridge_s0_translator:av_waitrequest
	wire    [0:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                        // peripheral_bridge_s0_translator:av_burstcount -> peripheral_bridge:s0_burstcount
	wire   [31:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata;                                         // peripheral_bridge_s0_translator:av_writedata -> peripheral_bridge:s0_writedata
	wire   [10:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_address;                                           // peripheral_bridge_s0_translator:av_address -> peripheral_bridge:s0_address
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_write;                                             // peripheral_bridge_s0_translator:av_write -> peripheral_bridge:s0_write
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_read;                                              // peripheral_bridge_s0_translator:av_read -> peripheral_bridge:s0_read
	wire   [31:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata;                                          // peripheral_bridge:s0_readdata -> peripheral_bridge_s0_translator:av_readdata
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                       // peripheral_bridge_s0_translator:av_debugaccess -> peripheral_bridge:s0_debugaccess
	wire          peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                     // peripheral_bridge:s0_readdatavalid -> peripheral_bridge_s0_translator:av_readdatavalid
	wire    [3:0] peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                        // peripheral_bridge_s0_translator:av_byteenable -> peripheral_bridge:s0_byteenable
	wire    [0:0] peripheral_bridge_m0_burstcount;                                                                       // peripheral_bridge:m0_burstcount -> peripheral_bridge_m0_translator:av_burstcount
	wire          peripheral_bridge_m0_waitrequest;                                                                      // peripheral_bridge_m0_translator:av_waitrequest -> peripheral_bridge:m0_waitrequest
	wire   [10:0] peripheral_bridge_m0_address;                                                                          // peripheral_bridge:m0_address -> peripheral_bridge_m0_translator:av_address
	wire   [31:0] peripheral_bridge_m0_writedata;                                                                        // peripheral_bridge:m0_writedata -> peripheral_bridge_m0_translator:av_writedata
	wire          peripheral_bridge_m0_write;                                                                            // peripheral_bridge:m0_write -> peripheral_bridge_m0_translator:av_write
	wire          peripheral_bridge_m0_read;                                                                             // peripheral_bridge:m0_read -> peripheral_bridge_m0_translator:av_read
	wire   [31:0] peripheral_bridge_m0_readdata;                                                                         // peripheral_bridge_m0_translator:av_readdata -> peripheral_bridge:m0_readdata
	wire          peripheral_bridge_m0_debugaccess;                                                                      // peripheral_bridge:m0_debugaccess -> peripheral_bridge_m0_translator:av_debugaccess
	wire    [3:0] peripheral_bridge_m0_byteenable;                                                                       // peripheral_bridge:m0_byteenable -> peripheral_bridge_m0_translator:av_byteenable
	wire          peripheral_bridge_m0_readdatavalid;                                                                    // peripheral_bridge_m0_translator:av_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire   [31:0] sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_writedata;                              // sd_card_controller_avalon_slave_translator:av_writedata -> sd_card_controller:avalon_slave_writedata
	wire    [7:0] sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_address;                                // sd_card_controller_avalon_slave_translator:av_address -> sd_card_controller:avalon_slave_address
	wire          sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_chipselect;                             // sd_card_controller_avalon_slave_translator:av_chipselect -> sd_card_controller:avalon_slave_chipselect
	wire          sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_write;                                  // sd_card_controller_avalon_slave_translator:av_write -> sd_card_controller:avalon_slave_write
	wire          sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_read;                                   // sd_card_controller_avalon_slave_translator:av_read -> sd_card_controller:avalon_slave_read
	wire   [31:0] sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_readdata;                               // sd_card_controller:avalon_slave_readdata -> sd_card_controller_avalon_slave_translator:av_readdata
	wire    [3:0] sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_byteenable;                             // sd_card_controller_avalon_slave_translator:av_byteenable -> sd_card_controller:avalon_slave_byteenable
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_anti_slave_0_writedata;                                               // lcd_i2c_scl_s1_translator:av_writedata -> lcd_i2c_scl:writedata
	wire    [1:0] lcd_i2c_scl_s1_translator_avalon_anti_slave_0_address;                                                 // lcd_i2c_scl_s1_translator:av_address -> lcd_i2c_scl:address
	wire          lcd_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect;                                              // lcd_i2c_scl_s1_translator:av_chipselect -> lcd_i2c_scl:chipselect
	wire          lcd_i2c_scl_s1_translator_avalon_anti_slave_0_write;                                                   // lcd_i2c_scl_s1_translator:av_write -> lcd_i2c_scl:write_n
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_anti_slave_0_readdata;                                                // lcd_i2c_scl:readdata -> lcd_i2c_scl_s1_translator:av_readdata
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_anti_slave_0_writedata;                                                // lcd_i2c_en_s1_translator:av_writedata -> lcd_i2c_en:writedata
	wire    [1:0] lcd_i2c_en_s1_translator_avalon_anti_slave_0_address;                                                  // lcd_i2c_en_s1_translator:av_address -> lcd_i2c_en:address
	wire          lcd_i2c_en_s1_translator_avalon_anti_slave_0_chipselect;                                               // lcd_i2c_en_s1_translator:av_chipselect -> lcd_i2c_en:chipselect
	wire          lcd_i2c_en_s1_translator_avalon_anti_slave_0_write;                                                    // lcd_i2c_en_s1_translator:av_write -> lcd_i2c_en:write_n
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_anti_slave_0_readdata;                                                 // lcd_i2c_en:readdata -> lcd_i2c_en_s1_translator:av_readdata
	wire   [31:0] lcd_i2c_sda_s1_translator_avalon_anti_slave_0_writedata;                                               // lcd_i2c_sda_s1_translator:av_writedata -> lcd_i2c_sda:writedata
	wire    [1:0] lcd_i2c_sda_s1_translator_avalon_anti_slave_0_address;                                                 // lcd_i2c_sda_s1_translator:av_address -> lcd_i2c_sda:address
	wire          lcd_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect;                                              // lcd_i2c_sda_s1_translator:av_chipselect -> lcd_i2c_sda:chipselect
	wire          lcd_i2c_sda_s1_translator_avalon_anti_slave_0_write;                                                   // lcd_i2c_sda_s1_translator:av_write -> lcd_i2c_sda:write_n
	wire   [31:0] lcd_i2c_sda_s1_translator_avalon_anti_slave_0_readdata;                                                // lcd_i2c_sda:readdata -> lcd_i2c_sda_s1_translator:av_readdata
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata;                                             // sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	wire    [2:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_address;                                               // sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect;                                            // sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_write;                                                 // sys_clk_timer_s1_translator:av_write -> sys_clk_timer:write_n
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata;                                              // sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	wire   [15:0] touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_writedata;                             // touch_panel_spi_spi_control_port_translator:av_writedata -> touch_panel_spi:data_from_cpu
	wire    [2:0] touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_address;                               // touch_panel_spi_spi_control_port_translator:av_address -> touch_panel_spi:mem_addr
	wire          touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_chipselect;                            // touch_panel_spi_spi_control_port_translator:av_chipselect -> touch_panel_spi:spi_select
	wire          touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_write;                                 // touch_panel_spi_spi_control_port_translator:av_write -> touch_panel_spi:write_n
	wire          touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_read;                                  // touch_panel_spi_spi_control_port_translator:av_read -> touch_panel_spi:read_n
	wire   [15:0] touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_readdata;                              // touch_panel_spi:data_to_cpu -> touch_panel_spi_spi_control_port_translator:av_readdata
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_writedata;                                     // touch_panel_pen_irq_n_s1_translator:av_writedata -> touch_panel_pen_irq_n:writedata
	wire    [1:0] touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_address;                                       // touch_panel_pen_irq_n_s1_translator:av_address -> touch_panel_pen_irq_n:address
	wire          touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_chipselect;                                    // touch_panel_pen_irq_n_s1_translator:av_chipselect -> touch_panel_pen_irq_n:chipselect
	wire          touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_write;                                         // touch_panel_pen_irq_n_s1_translator:av_write -> touch_panel_pen_irq_n:write_n
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_readdata;                                      // touch_panel_pen_irq_n:readdata -> touch_panel_pen_irq_n_s1_translator:av_readdata
	wire    [1:0] touch_panel_busy_s1_translator_avalon_anti_slave_0_address;                                            // touch_panel_busy_s1_translator:av_address -> touch_panel_busy:address
	wire   [31:0] touch_panel_busy_s1_translator_avalon_anti_slave_0_readdata;                                           // touch_panel_busy:readdata -> touch_panel_busy_s1_translator:av_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                               // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                 // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                   // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                      // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                     // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                      // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                  // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                               // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                      // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                       // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                        // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                          // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                             // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                            // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                             // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                         // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                      // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                       // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_waitrequest;                         // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_pixel_descriptor_write_translator:uav_waitrequest
	wire    [2:0] sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_burstcount;                          // sgdma_pixel_descriptor_write_translator:uav_burstcount -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_writedata;                           // sgdma_pixel_descriptor_write_translator:uav_writedata -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_address;                             // sgdma_pixel_descriptor_write_translator:uav_address -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_lock;                                // sgdma_pixel_descriptor_write_translator:uav_lock -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_write;                               // sgdma_pixel_descriptor_write_translator:uav_write -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_read;                                // sgdma_pixel_descriptor_write_translator:uav_read -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_readdata;                            // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_pixel_descriptor_write_translator:uav_readdata
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_debugaccess;                         // sgdma_pixel_descriptor_write_translator:uav_debugaccess -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_byteenable;                          // sgdma_pixel_descriptor_write_translator:uav_byteenable -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_readdatavalid;                       // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_pixel_descriptor_write_translator:uav_readdatavalid
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_waitrequest;                          // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_pixel_descriptor_read_translator:uav_waitrequest
	wire    [2:0] sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_burstcount;                           // sgdma_pixel_descriptor_read_translator:uav_burstcount -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_writedata;                            // sgdma_pixel_descriptor_read_translator:uav_writedata -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_address;                              // sgdma_pixel_descriptor_read_translator:uav_address -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_lock;                                 // sgdma_pixel_descriptor_read_translator:uav_lock -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_write;                                // sgdma_pixel_descriptor_read_translator:uav_write -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_read;                                 // sgdma_pixel_descriptor_read_translator:uav_read -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_readdata;                             // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_pixel_descriptor_read_translator:uav_readdata
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_debugaccess;                          // sgdma_pixel_descriptor_read_translator:uav_debugaccess -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_byteenable;                           // sgdma_pixel_descriptor_read_translator:uav_byteenable -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_readdatavalid;                        // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_pixel_descriptor_read_translator:uav_readdatavalid
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_waitrequest;                                   // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_pixel_m_read_translator:uav_waitrequest
	wire    [2:0] sgdma_pixel_m_read_translator_avalon_universal_master_0_burstcount;                                    // sgdma_pixel_m_read_translator:uav_burstcount -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] sgdma_pixel_m_read_translator_avalon_universal_master_0_writedata;                                     // sgdma_pixel_m_read_translator:uav_writedata -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] sgdma_pixel_m_read_translator_avalon_universal_master_0_address;                                       // sgdma_pixel_m_read_translator:uav_address -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_address
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_lock;                                          // sgdma_pixel_m_read_translator:uav_lock -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_lock
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_write;                                         // sgdma_pixel_m_read_translator:uav_write -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_write
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_read;                                          // sgdma_pixel_m_read_translator:uav_read -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] sgdma_pixel_m_read_translator_avalon_universal_master_0_readdata;                                      // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_pixel_m_read_translator:uav_readdata
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_debugaccess;                                   // sgdma_pixel_m_read_translator:uav_debugaccess -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] sgdma_pixel_m_read_translator_avalon_universal_master_0_byteenable;                                    // sgdma_pixel_m_read_translator:uav_byteenable -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_readdatavalid;                                 // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_pixel_m_read_translator:uav_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                           // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // sram_avalon_slave_translator:uav_waitrequest -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_avalon_slave_translator:uav_burstcount
	wire   [15:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                              // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_avalon_slave_translator:uav_writedata
	wire   [31:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> sram_avalon_slave_translator:uav_address
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                  // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> sram_avalon_slave_translator:uav_write
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                   // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sram_avalon_slave_translator:uav_lock
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                   // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> sram_avalon_slave_translator:uav_read
	wire   [15:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                               // sram_avalon_slave_translator:uav_readdata -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // sram_avalon_slave_translator:uav_readdatavalid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_avalon_slave_translator:uav_debugaccess
	wire    [1:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // sram_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_avalon_slave_translator:uav_byteenable
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                            // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [3:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // cfi_flash_uas_translator:uav_waitrequest -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_uas_translator:uav_burstcount
	wire    [7:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_uas_translator:uav_writedata
	wire   [31:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_address;                                    // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_uas_translator:uav_address
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_write;                                      // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_uas_translator:uav_write
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                       // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_uas_translator:uav_lock
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_read;                                       // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_uas_translator:uav_read
	wire    [7:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // cfi_flash_uas_translator:uav_readdata -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // cfi_flash_uas_translator:uav_readdatavalid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_uas_translator:uav_debugaccess
	wire    [0:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // cfi_flash_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_uas_translator:uav_byteenable
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [80:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [80:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire    [9:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // pll_pll_slave_translator:uav_waitrequest -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pll_pll_slave_translator:uav_burstcount
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pll_pll_slave_translator:uav_writedata
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                                    // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> pll_pll_slave_translator:uav_address
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                                      // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> pll_pll_slave_translator:uav_write
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pll_pll_slave_translator:uav_lock
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> pll_pll_slave_translator:uav_read
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // pll_pll_slave_translator:uav_readdata -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // pll_pll_slave_translator:uav_readdatavalid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pll_pll_slave_translator:uav_debugaccess
	wire    [3:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pll_pll_slave_translator:uav_byteenable
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                          // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                          // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // sgdma_pixel_csr_translator:uav_waitrequest -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_pixel_csr_translator:uav_burstcount
	wire   [31:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_pixel_csr_translator:uav_writedata
	wire   [31:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_address;                                  // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_pixel_csr_translator:uav_address
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_write;                                    // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_pixel_csr_translator:uav_write
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                     // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_pixel_csr_translator:uav_lock
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_read;                                     // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_pixel_csr_translator:uav_read
	wire   [31:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // sgdma_pixel_csr_translator:uav_readdata -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // sgdma_pixel_csr_translator:uav_readdatavalid -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_pixel_csr_translator:uav_debugaccess
	wire    [3:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_pixel_csr_translator:uav_byteenable
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                              // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // fifo_in_csr_translator:uav_waitrequest -> fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> fifo_in_csr_translator:uav_burstcount
	wire   [31:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> fifo_in_csr_translator:uav_writedata
	wire   [31:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_address;                                      // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_address -> fifo_in_csr_translator:uav_address
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_write;                                        // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_write -> fifo_in_csr_translator:uav_write
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_lock;                                         // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_lock -> fifo_in_csr_translator:uav_lock
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_read;                                         // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_read -> fifo_in_csr_translator:uav_read
	wire   [31:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // fifo_in_csr_translator:uav_readdata -> fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // fifo_in_csr_translator:uav_readdatavalid -> fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fifo_in_csr_translator:uav_debugaccess
	wire    [3:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // fifo_in_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> fifo_in_csr_translator:uav_byteenable
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // fifo_in_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                     // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                              // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                             // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // descriptor_mem_s1_translator:uav_waitrequest -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_mem_s1_translator:uav_burstcount
	wire   [31:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_mem_s1_translator:uav_writedata
	wire   [31:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_mem_s1_translator:uav_address
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_mem_s1_translator:uav_write
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_mem_s1_translator:uav_lock
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_mem_s1_translator:uav_read
	wire   [31:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // descriptor_mem_s1_translator:uav_readdata -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // descriptor_mem_s1_translator:uav_readdatavalid -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_mem_s1_translator:uav_debugaccess
	wire    [3:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_mem_s1_translator:uav_byteenable
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // peripheral_bridge_s0_translator:uav_waitrequest -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> peripheral_bridge_s0_translator:uav_burstcount
	wire   [31:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                           // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> peripheral_bridge_s0_translator:uav_writedata
	wire   [31:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                             // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> peripheral_bridge_s0_translator:uav_address
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                               // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> peripheral_bridge_s0_translator:uav_write
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                                // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> peripheral_bridge_s0_translator:uav_lock
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                                // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> peripheral_bridge_s0_translator:uav_read
	wire   [31:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                            // peripheral_bridge_s0_translator:uav_readdata -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // peripheral_bridge_s0_translator:uav_readdatavalid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> peripheral_bridge_s0_translator:uav_debugaccess
	wire    [3:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> peripheral_bridge_s0_translator:uav_byteenable
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                         // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest;                                 // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> peripheral_bridge_m0_translator:uav_waitrequest
	wire    [2:0] peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount;                                  // peripheral_bridge_m0_translator:uav_burstcount -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] peripheral_bridge_m0_translator_avalon_universal_master_0_writedata;                                   // peripheral_bridge_m0_translator:uav_writedata -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [10:0] peripheral_bridge_m0_translator_avalon_universal_master_0_address;                                     // peripheral_bridge_m0_translator:uav_address -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_lock;                                        // peripheral_bridge_m0_translator:uav_lock -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_write;                                       // peripheral_bridge_m0_translator:uav_write -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_read;                                        // peripheral_bridge_m0_translator:uav_read -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] peripheral_bridge_m0_translator_avalon_universal_master_0_readdata;                                    // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> peripheral_bridge_m0_translator:uav_readdata
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess;                                 // peripheral_bridge_m0_translator:uav_debugaccess -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable;                                  // peripheral_bridge_m0_translator:uav_byteenable -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                               // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> peripheral_bridge_m0_translator:uav_readdatavalid
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // sd_card_controller_avalon_slave_translator:uav_waitrequest -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sd_card_controller_avalon_slave_translator:uav_burstcount
	wire   [31:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sd_card_controller_avalon_slave_translator:uav_writedata
	wire   [10:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> sd_card_controller_avalon_slave_translator:uav_address
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> sd_card_controller_avalon_slave_translator:uav_write
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sd_card_controller_avalon_slave_translator:uav_lock
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> sd_card_controller_avalon_slave_translator:uav_read
	wire   [31:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // sd_card_controller_avalon_slave_translator:uav_readdata -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // sd_card_controller_avalon_slave_translator:uav_readdatavalid -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sd_card_controller_avalon_slave_translator:uav_debugaccess
	wire    [3:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sd_card_controller_avalon_slave_translator:uav_byteenable
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // lcd_i2c_scl_s1_translator:uav_waitrequest -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_i2c_scl_s1_translator:uav_burstcount
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_i2c_scl_s1_translator:uav_writedata
	wire   [10:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_i2c_scl_s1_translator:uav_address
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_i2c_scl_s1_translator:uav_write
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_i2c_scl_s1_translator:uav_lock
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_i2c_scl_s1_translator:uav_read
	wire   [31:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // lcd_i2c_scl_s1_translator:uav_readdata -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // lcd_i2c_scl_s1_translator:uav_readdatavalid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_i2c_scl_s1_translator:uav_debugaccess
	wire    [3:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_i2c_scl_s1_translator:uav_byteenable
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // lcd_i2c_en_s1_translator:uav_waitrequest -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_i2c_en_s1_translator:uav_burstcount
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_i2c_en_s1_translator:uav_writedata
	wire   [10:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_i2c_en_s1_translator:uav_address
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_i2c_en_s1_translator:uav_write
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_i2c_en_s1_translator:uav_lock
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_i2c_en_s1_translator:uav_read
	wire   [31:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // lcd_i2c_en_s1_translator:uav_readdata -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // lcd_i2c_en_s1_translator:uav_readdatavalid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_i2c_en_s1_translator:uav_debugaccess
	wire    [3:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_i2c_en_s1_translator:uav_byteenable
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // lcd_i2c_sda_s1_translator:uav_waitrequest -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_i2c_sda_s1_translator:uav_burstcount
	wire   [31:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_i2c_sda_s1_translator:uav_writedata
	wire   [10:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_address -> lcd_i2c_sda_s1_translator:uav_address
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_write -> lcd_i2c_sda_s1_translator:uav_write
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_i2c_sda_s1_translator:uav_lock
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_read -> lcd_i2c_sda_s1_translator:uav_read
	wire   [31:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // lcd_i2c_sda_s1_translator:uav_readdata -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // lcd_i2c_sda_s1_translator:uav_readdatavalid -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_i2c_sda_s1_translator:uav_debugaccess
	wire    [3:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_i2c_sda_s1_translator:uav_byteenable
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	wire   [10:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	wire    [3:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // touch_panel_spi_spi_control_port_translator:uav_waitrequest -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> touch_panel_spi_spi_control_port_translator:uav_burstcount
	wire   [31:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> touch_panel_spi_spi_control_port_translator:uav_writedata
	wire   [10:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_address -> touch_panel_spi_spi_control_port_translator:uav_address
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_write -> touch_panel_spi_spi_control_port_translator:uav_write
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> touch_panel_spi_spi_control_port_translator:uav_lock
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_read -> touch_panel_spi_spi_control_port_translator:uav_read
	wire   [31:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // touch_panel_spi_spi_control_port_translator:uav_readdata -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // touch_panel_spi_spi_control_port_translator:uav_readdatavalid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> touch_panel_spi_spi_control_port_translator:uav_debugaccess
	wire    [3:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> touch_panel_spi_spi_control_port_translator:uav_byteenable
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // touch_panel_pen_irq_n_s1_translator:uav_waitrequest -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> touch_panel_pen_irq_n_s1_translator:uav_burstcount
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> touch_panel_pen_irq_n_s1_translator:uav_writedata
	wire   [10:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_address -> touch_panel_pen_irq_n_s1_translator:uav_address
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_write -> touch_panel_pen_irq_n_s1_translator:uav_write
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_lock -> touch_panel_pen_irq_n_s1_translator:uav_lock
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_read -> touch_panel_pen_irq_n_s1_translator:uav_read
	wire   [31:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // touch_panel_pen_irq_n_s1_translator:uav_readdata -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // touch_panel_pen_irq_n_s1_translator:uav_readdatavalid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> touch_panel_pen_irq_n_s1_translator:uav_debugaccess
	wire    [3:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> touch_panel_pen_irq_n_s1_translator:uav_byteenable
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // touch_panel_busy_s1_translator:uav_waitrequest -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> touch_panel_busy_s1_translator:uav_burstcount
	wire   [31:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> touch_panel_busy_s1_translator:uav_writedata
	wire   [10:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_address -> touch_panel_busy_s1_translator:uav_address
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_write -> touch_panel_busy_s1_translator:uav_write
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_lock -> touch_panel_busy_s1_translator:uav_lock
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_read -> touch_panel_busy_s1_translator:uav_read
	wire   [31:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // touch_panel_busy_s1_translator:uav_readdata -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // touch_panel_busy_s1_translator:uav_readdatavalid -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> touch_panel_busy_s1_translator:uav_debugaccess
	wire    [3:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> touch_panel_busy_s1_translator:uav_byteenable
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                            // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [106:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                             // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                   // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                           // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [106:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                   // addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket;                // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid;                      // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket;              // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [106:0] sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_data;                       // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router_002:sink_ready -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                 // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid;                       // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket;               // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [106:0] sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_data;                        // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready;                       // addr_router_003:sink_ready -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket;                          // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_valid;                                // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket;                        // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [106:0] sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_data;                                 // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_ready;                                // addr_router_004:sink_ready -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                              // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [106:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                  // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [88:0] sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                   // sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_001:sink_ready -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                           // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [106:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                            // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                      // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [79:0] cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_data;                                       // cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_003:sink_ready -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                      // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [106:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_004:sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                    // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [106:0] sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_data;                                     // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_005:sink_ready -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_valid;                                        // fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_data;                                         // fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_006:sink_ready -> fifo_in_csr_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [106:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router_007:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [106:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_008:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [106:0] descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_009:sink_ready -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                               // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [106:0] peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                                // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_010:sink_ready -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                        // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                              // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                      // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire   [81:0] peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                               // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                              // addr_router_005:sink_ready -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [81:0] sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_011:sink_ready -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire   [81:0] lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_012:sink_ready -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [81:0] lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_013:sink_ready -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [81:0] lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_014:sink_ready -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [81:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_015:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [81:0] touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_016:sink_ready -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire   [81:0] touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_017:sink_ready -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire   [81:0] touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_018:sink_ready -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                           // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                 // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                         // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [106:0] addr_router_src_data;                                                                                  // addr_router:src_data -> limiter:cmd_sink_data
	wire   [10:0] addr_router_src_channel;                                                                               // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                 // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                           // limiter:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                 // limiter:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                         // limiter:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_rsp_src_data;                                                                                  // limiter:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] limiter_rsp_src_channel;                                                                               // limiter:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                 // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                       // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                             // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                     // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [106:0] addr_router_001_src_data;                                                                              // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [10:0] addr_router_001_src_channel;                                                                           // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                             // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                       // limiter_001:rsp_src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                             // limiter_001:rsp_src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                     // limiter_001:rsp_src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_001_rsp_src_data;                                                                              // limiter_001:rsp_src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] limiter_001_rsp_src_channel;                                                                           // limiter_001:rsp_src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                             // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_005_src_endofpacket;                                                                       // addr_router_005:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_005_src_valid;                                                                             // addr_router_005:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_005_src_startofpacket;                                                                     // addr_router_005:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire   [81:0] addr_router_005_src_data;                                                                              // addr_router_005:src_data -> limiter_002:cmd_sink_data
	wire    [7:0] addr_router_005_src_channel;                                                                           // addr_router_005:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_005_src_ready;                                                                             // limiter_002:cmd_sink_ready -> addr_router_005:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                       // limiter_002:rsp_src_endofpacket -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                             // limiter_002:rsp_src_valid -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                     // limiter_002:rsp_src_startofpacket -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [81:0] limiter_002_rsp_src_data;                                                                              // limiter_002:rsp_src_data -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [7:0] limiter_002_rsp_src_channel;                                                                           // limiter_002:rsp_src_channel -> peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                             // peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                     // burst_adapter:source0_endofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                           // burst_adapter:source0_valid -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                   // burst_adapter:source0_startofpacket -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_source0_data;                                                                            // burst_adapter:source0_data -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                           // sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [10:0] burst_adapter_source0_channel;                                                                         // burst_adapter:source0_channel -> sram_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                 // burst_adapter_001:source0_endofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                       // burst_adapter_001:source0_valid -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                               // burst_adapter_001:source0_startofpacket -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [79:0] burst_adapter_001_source0_data;                                                                        // burst_adapter_001:source0_data -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                       // cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [10:0] burst_adapter_001_source0_channel;                                                                     // burst_adapter_001:source0_channel -> cfi_flash_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                        // rst_controller:reset_out -> [crosser:out_reset, crosser_001:in_reset, id_router_004:reset, pll:reset, pll_pll_slave_translator:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_004:reset]
	wire          cpu_jtag_debug_module_reset_reset;                                                                     // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                                                    // rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, burst_adapter:reset, burst_adapter_001:reset, cfi_flash:reset_reset, cfi_flash_uas_translator:reset, cfi_flash_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_009:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:in_reset, crosser_001:out_reset, descriptor_mem:reset, descriptor_mem_s1_translator:reset, descriptor_mem_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fifo:wrreset_n, fifo_in_csr_translator:reset, fifo_in_csr_translator_avalon_universal_slave_0_agent:reset, fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, peripheral_bridge:s0_reset, peripheral_bridge_s0_translator:reset, peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:reset, peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_pixel:system_reset_n, sgdma_pixel_csr_translator:reset, sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_pixel_descriptor_read_translator:reset, sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_pixel_descriptor_write_translator:reset, sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_pixel_m_read_translator:reset, sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:reset, sram:reset_n, sram_avalon_slave_translator:reset, sram_avalon_slave_translator_avalon_universal_slave_0_agent:reset, sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timing_adapter:reset_n, tri_state_bridge_flash_bridge_0:reset, tri_state_bridge_flash_pinSharer_0:reset_reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_001_reset_out_reset_req;                                                                // rst_controller_001:reset_req -> descriptor_mem:reset_req
	wire          rst_controller_002_reset_out_reset;                                                                    // rst_controller_002:reset_out -> [fifo:rdreset_n, fifo_to_pixel_converter:reset_n, pixel_converter:reset_n, video_sync_generator:reset_n]
	wire          rst_controller_003_reset_out_reset;                                                                    // rst_controller_003:reset_out -> [addr_router_005:reset, cmd_xbar_demux_005:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, lcd_i2c_en:reset_n, lcd_i2c_en_s1_translator:reset, lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:reset, lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_i2c_scl:reset_n, lcd_i2c_scl_s1_translator:reset, lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:reset, lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_i2c_sda:reset_n, lcd_i2c_sda_s1_translator:reset, lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:reset, lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_002:reset, peripheral_bridge:m0_reset, peripheral_bridge_m0_translator:reset, peripheral_bridge_m0_translator_avalon_universal_master_0_agent:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_mux_005:reset, sd_card_controller:reset_n, sd_card_controller_avalon_slave_translator:reset, sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:reset, sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sys_clk_timer:reset_n, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, touch_panel_busy:reset_n, touch_panel_busy_s1_translator:reset, touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:reset, touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, touch_panel_pen_irq_n:reset_n, touch_panel_pen_irq_n_s1_translator:reset, touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:reset, touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, touch_panel_spi:reset_n, touch_panel_spi_spi_control_port_translator:reset, touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:reset, touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                       // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                             // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                     // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src0_data;                                                                              // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [10:0] cmd_xbar_demux_src0_channel;                                                                           // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                             // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                       // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                             // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                     // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src1_data;                                                                              // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [10:0] cmd_xbar_demux_src1_channel;                                                                           // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src1_ready;                                                                             // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                       // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                             // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                     // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src2_data;                                                                              // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [10:0] cmd_xbar_demux_src2_channel;                                                                           // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                             // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                       // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                             // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                     // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src3_data;                                                                              // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [10:0] cmd_xbar_demux_src3_channel;                                                                           // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                             // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                   // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                         // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                 // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src0_data;                                                                          // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [10:0] cmd_xbar_demux_001_src0_channel;                                                                       // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                         // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                   // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                         // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                 // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src1_data;                                                                          // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [10:0] cmd_xbar_demux_001_src1_channel;                                                                       // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                         // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                   // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                         // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                 // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src2_data;                                                                          // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [10:0] cmd_xbar_demux_001_src2_channel;                                                                       // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                         // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                   // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                         // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                 // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src3_data;                                                                          // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [10:0] cmd_xbar_demux_001_src3_channel;                                                                       // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                         // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                   // cmd_xbar_demux_001:src5_endofpacket -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                         // cmd_xbar_demux_001:src5_valid -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                 // cmd_xbar_demux_001:src5_startofpacket -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src5_data;                                                                          // cmd_xbar_demux_001:src5_data -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src5_channel;                                                                       // cmd_xbar_demux_001:src5_channel -> sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                   // cmd_xbar_demux_001:src6_endofpacket -> fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                         // cmd_xbar_demux_001:src6_valid -> fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                 // cmd_xbar_demux_001:src6_startofpacket -> fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src6_data;                                                                          // cmd_xbar_demux_001:src6_data -> fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src6_channel;                                                                       // cmd_xbar_demux_001:src6_channel -> fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                   // cmd_xbar_demux_001:src7_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                         // cmd_xbar_demux_001:src7_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                 // cmd_xbar_demux_001:src7_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src7_data;                                                                          // cmd_xbar_demux_001:src7_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src7_channel;                                                                       // cmd_xbar_demux_001:src7_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                   // cmd_xbar_demux_001:src8_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                         // cmd_xbar_demux_001:src8_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                 // cmd_xbar_demux_001:src8_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src8_data;                                                                          // cmd_xbar_demux_001:src8_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src8_channel;                                                                       // cmd_xbar_demux_001:src8_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                   // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                         // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                 // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src9_data;                                                                          // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink0_data
	wire   [10:0] cmd_xbar_demux_001_src9_channel;                                                                       // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire          cmd_xbar_demux_001_src9_ready;                                                                         // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux_001:src9_ready
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                  // cmd_xbar_demux_001:src10_endofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                        // cmd_xbar_demux_001:src10_valid -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                // cmd_xbar_demux_001:src10_startofpacket -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src10_data;                                                                         // cmd_xbar_demux_001:src10_data -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_001_src10_channel;                                                                      // cmd_xbar_demux_001:src10_channel -> peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                   // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                         // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_009:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                 // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src0_data;                                                                          // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_009:sink1_data
	wire   [10:0] cmd_xbar_demux_002_src0_channel;                                                                       // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_009:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                         // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                   // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_009:sink2_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                         // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_009:sink2_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                 // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_009:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src0_data;                                                                          // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_009:sink2_data
	wire   [10:0] cmd_xbar_demux_003_src0_channel;                                                                       // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_009:sink2_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                         // cmd_xbar_mux_009:sink2_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                   // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                         // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_002:sink2_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                 // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src0_data;                                                                          // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_002:sink2_data
	wire   [10:0] cmd_xbar_demux_004_src0_channel;                                                                       // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_002:sink2_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                         // cmd_xbar_mux_002:sink2_ready -> cmd_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                       // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                             // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                     // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src0_data;                                                                              // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [10:0] rsp_xbar_demux_src0_channel;                                                                           // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                             // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                       // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                             // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                     // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src1_data;                                                                              // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [10:0] rsp_xbar_demux_src1_channel;                                                                           // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                             // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                   // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                         // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                 // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src0_data;                                                                          // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [10:0] rsp_xbar_demux_001_src0_channel;                                                                       // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                         // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                   // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                         // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                 // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src1_data;                                                                          // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [10:0] rsp_xbar_demux_001_src1_channel;                                                                       // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                         // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                   // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                         // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                 // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src0_data;                                                                          // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [10:0] rsp_xbar_demux_002_src0_channel;                                                                       // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                         // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                   // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                         // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                 // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src1_data;                                                                          // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [10:0] rsp_xbar_demux_002_src1_channel;                                                                       // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                         // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_002_src2_endofpacket;                                                                   // rsp_xbar_demux_002:src2_endofpacket -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_002_src2_valid;                                                                         // rsp_xbar_demux_002:src2_valid -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_002_src2_startofpacket;                                                                 // rsp_xbar_demux_002:src2_startofpacket -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src2_data;                                                                          // rsp_xbar_demux_002:src2_data -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] rsp_xbar_demux_002_src2_channel;                                                                       // rsp_xbar_demux_002:src2_channel -> sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                   // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                         // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                 // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src0_data;                                                                          // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [10:0] rsp_xbar_demux_003_src0_channel;                                                                       // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                         // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                   // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                         // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                 // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src1_data;                                                                          // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [10:0] rsp_xbar_demux_003_src1_channel;                                                                       // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                         // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                   // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                         // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                 // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src0_data;                                                                          // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [10:0] rsp_xbar_demux_005_src0_channel;                                                                       // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                         // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                   // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                         // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                 // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                          // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire   [10:0] rsp_xbar_demux_006_src0_channel;                                                                       // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                         // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                   // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                         // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                 // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_007_src0_data;                                                                          // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [10:0] rsp_xbar_demux_007_src0_channel;                                                                       // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                         // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                   // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                         // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                 // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_008_src0_data;                                                                          // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [10:0] rsp_xbar_demux_008_src0_channel;                                                                       // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                         // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                   // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                         // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                 // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src0_data;                                                                          // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [10:0] rsp_xbar_demux_009_src0_channel;                                                                       // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                         // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_009_src1_endofpacket;                                                                   // rsp_xbar_demux_009:src1_endofpacket -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_009_src1_valid;                                                                         // rsp_xbar_demux_009:src1_valid -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_009_src1_startofpacket;                                                                 // rsp_xbar_demux_009:src1_startofpacket -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src1_data;                                                                          // rsp_xbar_demux_009:src1_data -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] rsp_xbar_demux_009_src1_channel;                                                                       // rsp_xbar_demux_009:src1_channel -> sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_009_src2_endofpacket;                                                                   // rsp_xbar_demux_009:src2_endofpacket -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_009_src2_valid;                                                                         // rsp_xbar_demux_009:src2_valid -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_009_src2_startofpacket;                                                                 // rsp_xbar_demux_009:src2_startofpacket -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src2_data;                                                                          // rsp_xbar_demux_009:src2_data -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] rsp_xbar_demux_009_src2_channel;                                                                       // rsp_xbar_demux_009:src2_channel -> sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                   // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                         // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                 // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src0_data;                                                                          // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [10:0] rsp_xbar_demux_010_src0_channel;                                                                       // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                         // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                           // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                         // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [106:0] limiter_cmd_src_data;                                                                                  // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [10:0] limiter_cmd_src_channel;                                                                               // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                 // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                          // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                        // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_src_data;                                                                                 // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [10:0] rsp_xbar_mux_src_channel;                                                                              // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                       // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                     // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [106:0] limiter_001_cmd_src_data;                                                                              // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [10:0] limiter_001_cmd_src_channel;                                                                           // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                             // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                      // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                            // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                    // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_001_src_data;                                                                             // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [10:0] rsp_xbar_mux_001_src_channel;                                                                          // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                            // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                       // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                             // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                     // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [106:0] addr_router_002_src_data;                                                                              // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [10:0] addr_router_002_src_channel;                                                                           // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                             // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_demux_009_src1_ready;                                                                         // sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_009:src1_ready
	wire          addr_router_003_src_endofpacket;                                                                       // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                             // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                     // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [106:0] addr_router_003_src_data;                                                                              // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [10:0] addr_router_003_src_channel;                                                                           // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                             // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_009_src2_ready;                                                                         // sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_009:src2_ready
	wire          addr_router_004_src_endofpacket;                                                                       // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                             // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                     // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [106:0] addr_router_004_src_data;                                                                              // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [10:0] addr_router_004_src_channel;                                                                           // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                             // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_002_src2_ready;                                                                         // sgdma_pixel_m_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_002:src2_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                          // cmd_xbar_mux:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                // cmd_xbar_mux:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                        // cmd_xbar_mux:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_src_data;                                                                                 // cmd_xbar_mux:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_mux_src_channel;                                                                              // cmd_xbar_mux:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                             // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                   // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                           // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [106:0] id_router_src_data;                                                                                    // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [10:0] id_router_src_channel;                                                                                 // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                   // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                      // cmd_xbar_mux_002:src_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                            // cmd_xbar_mux_002:src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                    // cmd_xbar_mux_002:src_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_002_src_data;                                                                             // cmd_xbar_mux_002:src_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_mux_002_src_channel;                                                                          // cmd_xbar_mux_002:src_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                            // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                         // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                               // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                       // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [106:0] id_router_002_src_data;                                                                                // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [10:0] id_router_002_src_channel;                                                                             // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                               // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          crosser_out_ready;                                                                                     // pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_004_src_endofpacket;                                                                         // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                               // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                       // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] id_router_004_src_data;                                                                                // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [10:0] id_router_004_src_channel;                                                                             // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                               // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                         // sgdma_pixel_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                         // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                               // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                       // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [106:0] id_router_005_src_data;                                                                                // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [10:0] id_router_005_src_channel;                                                                             // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                               // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_001_src6_ready;                                                                         // fifo_in_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire          id_router_006_src_endofpacket;                                                                         // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                               // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                       // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                                // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [10:0] id_router_006_src_channel;                                                                             // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                               // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                         // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                               // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                       // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [106:0] id_router_007_src_data;                                                                                // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [10:0] id_router_007_src_channel;                                                                             // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                               // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                         // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                               // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                       // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [106:0] id_router_008_src_data;                                                                                // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [10:0] id_router_008_src_channel;                                                                             // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                               // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_009_src_endofpacket;                                                                      // cmd_xbar_mux_009:src_endofpacket -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_009_src_valid;                                                                            // cmd_xbar_mux_009:src_valid -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_009_src_startofpacket;                                                                    // cmd_xbar_mux_009:src_startofpacket -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_009_src_data;                                                                             // cmd_xbar_mux_009:src_data -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_mux_009_src_channel;                                                                          // cmd_xbar_mux_009:src_channel -> descriptor_mem_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_009_src_ready;                                                                            // descriptor_mem_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire          id_router_009_src_endofpacket;                                                                         // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                               // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                       // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [106:0] id_router_009_src_data;                                                                                // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [10:0] id_router_009_src_channel;                                                                             // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                               // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_001_src10_ready;                                                                        // peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire          id_router_010_src_endofpacket;                                                                         // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                               // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                       // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [106:0] id_router_010_src_data;                                                                                // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [10:0] id_router_010_src_channel;                                                                             // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                               // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                   // cmd_xbar_demux_005:src0_endofpacket -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                         // cmd_xbar_demux_005:src0_valid -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                 // cmd_xbar_demux_005:src0_startofpacket -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src0_data;                                                                          // cmd_xbar_demux_005:src0_data -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src0_channel;                                                                       // cmd_xbar_demux_005:src0_channel -> sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src1_endofpacket;                                                                   // cmd_xbar_demux_005:src1_endofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src1_valid;                                                                         // cmd_xbar_demux_005:src1_valid -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src1_startofpacket;                                                                 // cmd_xbar_demux_005:src1_startofpacket -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src1_data;                                                                          // cmd_xbar_demux_005:src1_data -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src1_channel;                                                                       // cmd_xbar_demux_005:src1_channel -> lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src2_endofpacket;                                                                   // cmd_xbar_demux_005:src2_endofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src2_valid;                                                                         // cmd_xbar_demux_005:src2_valid -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src2_startofpacket;                                                                 // cmd_xbar_demux_005:src2_startofpacket -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src2_data;                                                                          // cmd_xbar_demux_005:src2_data -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src2_channel;                                                                       // cmd_xbar_demux_005:src2_channel -> lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src3_endofpacket;                                                                   // cmd_xbar_demux_005:src3_endofpacket -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src3_valid;                                                                         // cmd_xbar_demux_005:src3_valid -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src3_startofpacket;                                                                 // cmd_xbar_demux_005:src3_startofpacket -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src3_data;                                                                          // cmd_xbar_demux_005:src3_data -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src3_channel;                                                                       // cmd_xbar_demux_005:src3_channel -> lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src4_endofpacket;                                                                   // cmd_xbar_demux_005:src4_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src4_valid;                                                                         // cmd_xbar_demux_005:src4_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src4_startofpacket;                                                                 // cmd_xbar_demux_005:src4_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src4_data;                                                                          // cmd_xbar_demux_005:src4_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src4_channel;                                                                       // cmd_xbar_demux_005:src4_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src5_endofpacket;                                                                   // cmd_xbar_demux_005:src5_endofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src5_valid;                                                                         // cmd_xbar_demux_005:src5_valid -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src5_startofpacket;                                                                 // cmd_xbar_demux_005:src5_startofpacket -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src5_data;                                                                          // cmd_xbar_demux_005:src5_data -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src5_channel;                                                                       // cmd_xbar_demux_005:src5_channel -> touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src6_endofpacket;                                                                   // cmd_xbar_demux_005:src6_endofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src6_valid;                                                                         // cmd_xbar_demux_005:src6_valid -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src6_startofpacket;                                                                 // cmd_xbar_demux_005:src6_startofpacket -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src6_data;                                                                          // cmd_xbar_demux_005:src6_data -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src6_channel;                                                                       // cmd_xbar_demux_005:src6_channel -> touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_005_src7_endofpacket;                                                                   // cmd_xbar_demux_005:src7_endofpacket -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_005_src7_valid;                                                                         // cmd_xbar_demux_005:src7_valid -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_005_src7_startofpacket;                                                                 // cmd_xbar_demux_005:src7_startofpacket -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] cmd_xbar_demux_005_src7_data;                                                                          // cmd_xbar_demux_005:src7_data -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [7:0] cmd_xbar_demux_005_src7_channel;                                                                       // cmd_xbar_demux_005:src7_channel -> touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                   // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_005:sink0_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                         // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_005:sink0_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                 // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_005:sink0_startofpacket
	wire   [81:0] rsp_xbar_demux_011_src0_data;                                                                          // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_005:sink0_data
	wire    [7:0] rsp_xbar_demux_011_src0_channel;                                                                       // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_005:sink0_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                         // rsp_xbar_mux_005:sink0_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                   // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_005:sink1_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                         // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_005:sink1_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                 // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_005:sink1_startofpacket
	wire   [81:0] rsp_xbar_demux_012_src0_data;                                                                          // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_005:sink1_data
	wire    [7:0] rsp_xbar_demux_012_src0_channel;                                                                       // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_005:sink1_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                         // rsp_xbar_mux_005:sink1_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                   // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_005:sink2_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                         // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_005:sink2_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                 // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_005:sink2_startofpacket
	wire   [81:0] rsp_xbar_demux_013_src0_data;                                                                          // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_005:sink2_data
	wire    [7:0] rsp_xbar_demux_013_src0_channel;                                                                       // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_005:sink2_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                         // rsp_xbar_mux_005:sink2_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                   // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_005:sink3_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                         // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_005:sink3_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                 // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_005:sink3_startofpacket
	wire   [81:0] rsp_xbar_demux_014_src0_data;                                                                          // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_005:sink3_data
	wire    [7:0] rsp_xbar_demux_014_src0_channel;                                                                       // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_005:sink3_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                         // rsp_xbar_mux_005:sink3_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                   // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_005:sink4_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                         // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_005:sink4_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                 // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_005:sink4_startofpacket
	wire   [81:0] rsp_xbar_demux_015_src0_data;                                                                          // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_005:sink4_data
	wire    [7:0] rsp_xbar_demux_015_src0_channel;                                                                       // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_005:sink4_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                         // rsp_xbar_mux_005:sink4_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                   // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_005:sink5_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                         // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_005:sink5_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                 // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_005:sink5_startofpacket
	wire   [81:0] rsp_xbar_demux_016_src0_data;                                                                          // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_005:sink5_data
	wire    [7:0] rsp_xbar_demux_016_src0_channel;                                                                       // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_005:sink5_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                         // rsp_xbar_mux_005:sink5_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                   // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_005:sink6_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                         // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_005:sink6_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                 // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_005:sink6_startofpacket
	wire   [81:0] rsp_xbar_demux_017_src0_data;                                                                          // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_005:sink6_data
	wire    [7:0] rsp_xbar_demux_017_src0_channel;                                                                       // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_005:sink6_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                         // rsp_xbar_mux_005:sink6_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                   // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_005:sink7_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                         // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_005:sink7_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                 // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_005:sink7_startofpacket
	wire   [81:0] rsp_xbar_demux_018_src0_data;                                                                          // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_005:sink7_data
	wire    [7:0] rsp_xbar_demux_018_src0_channel;                                                                       // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_005:sink7_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                         // rsp_xbar_mux_005:sink7_ready -> rsp_xbar_demux_018:src0_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                       // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                     // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire   [81:0] limiter_002_cmd_src_data;                                                                              // limiter_002:cmd_src_data -> cmd_xbar_demux_005:sink_data
	wire    [7:0] limiter_002_cmd_src_channel;                                                                           // limiter_002:cmd_src_channel -> cmd_xbar_demux_005:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                             // cmd_xbar_demux_005:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_005_src_endofpacket;                                                                      // rsp_xbar_mux_005:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_005_src_valid;                                                                            // rsp_xbar_mux_005:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_005_src_startofpacket;                                                                    // rsp_xbar_mux_005:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire   [81:0] rsp_xbar_mux_005_src_data;                                                                             // rsp_xbar_mux_005:src_data -> limiter_002:rsp_sink_data
	wire    [7:0] rsp_xbar_mux_005_src_channel;                                                                          // rsp_xbar_mux_005:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_005_src_ready;                                                                            // limiter_002:rsp_sink_ready -> rsp_xbar_mux_005:src_ready
	wire          cmd_xbar_demux_005_src0_ready;                                                                         // sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src0_ready
	wire          id_router_011_src_endofpacket;                                                                         // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                               // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                       // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [81:0] id_router_011_src_data;                                                                                // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire    [7:0] id_router_011_src_channel;                                                                             // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                               // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_005_src1_ready;                                                                         // lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src1_ready
	wire          id_router_012_src_endofpacket;                                                                         // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                               // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                       // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [81:0] id_router_012_src_data;                                                                                // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire    [7:0] id_router_012_src_channel;                                                                             // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                               // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_005_src2_ready;                                                                         // lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src2_ready
	wire          id_router_013_src_endofpacket;                                                                         // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                               // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                       // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [81:0] id_router_013_src_data;                                                                                // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire    [7:0] id_router_013_src_channel;                                                                             // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                               // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_005_src3_ready;                                                                         // lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src3_ready
	wire          id_router_014_src_endofpacket;                                                                         // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                               // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                       // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [81:0] id_router_014_src_data;                                                                                // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire    [7:0] id_router_014_src_channel;                                                                             // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                               // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_005_src4_ready;                                                                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src4_ready
	wire          id_router_015_src_endofpacket;                                                                         // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                               // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                       // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [81:0] id_router_015_src_data;                                                                                // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire    [7:0] id_router_015_src_channel;                                                                             // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                               // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_005_src5_ready;                                                                         // touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src5_ready
	wire          id_router_016_src_endofpacket;                                                                         // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                               // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                       // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire   [81:0] id_router_016_src_data;                                                                                // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire    [7:0] id_router_016_src_channel;                                                                             // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                               // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_005_src6_ready;                                                                         // touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src6_ready
	wire          id_router_017_src_endofpacket;                                                                         // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                               // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                       // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire   [81:0] id_router_017_src_data;                                                                                // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire    [7:0] id_router_017_src_channel;                                                                             // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                               // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_005_src7_ready;                                                                         // touch_panel_busy_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_005:src7_ready
	wire          id_router_018_src_endofpacket;                                                                         // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                               // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                       // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire   [81:0] id_router_018_src_data;                                                                                // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire    [7:0] id_router_018_src_channel;                                                                             // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                               // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                      // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                            // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                    // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [106:0] cmd_xbar_mux_001_src_data;                                                                             // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire   [10:0] cmd_xbar_mux_001_src_channel;                                                                          // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                            // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire          width_adapter_src_endofpacket;                                                                         // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                               // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                       // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [88:0] width_adapter_src_data;                                                                                // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                               // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [10:0] width_adapter_src_channel;                                                                             // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_001_src_endofpacket;                                                                         // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_001_src_valid;                                                                               // id_router_001:src_valid -> width_adapter_001:in_valid
	wire          id_router_001_src_startofpacket;                                                                       // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire   [88:0] id_router_001_src_data;                                                                                // id_router_001:src_data -> width_adapter_001:in_data
	wire   [10:0] id_router_001_src_channel;                                                                             // id_router_001:src_channel -> width_adapter_001:in_channel
	wire          id_router_001_src_ready;                                                                               // width_adapter_001:in_ready -> id_router_001:src_ready
	wire          width_adapter_001_src_endofpacket;                                                                     // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                                           // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                                   // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [106:0] width_adapter_001_src_data;                                                                            // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_001_src_ready;                                                                           // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [10:0] width_adapter_001_src_channel;                                                                         // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                      // cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                            // cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                    // cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [106:0] cmd_xbar_mux_003_src_data;                                                                             // cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	wire   [10:0] cmd_xbar_mux_003_src_channel;                                                                          // cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                            // width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	wire          width_adapter_002_src_endofpacket;                                                                     // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                           // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                   // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [79:0] width_adapter_002_src_data;                                                                            // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                                           // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire   [10:0] width_adapter_002_src_channel;                                                                         // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_003_src_endofpacket;                                                                         // id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_003_src_valid;                                                                               // id_router_003:src_valid -> width_adapter_003:in_valid
	wire          id_router_003_src_startofpacket;                                                                       // id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	wire   [79:0] id_router_003_src_data;                                                                                // id_router_003:src_data -> width_adapter_003:in_data
	wire   [10:0] id_router_003_src_channel;                                                                             // id_router_003:src_channel -> width_adapter_003:in_channel
	wire          id_router_003_src_ready;                                                                               // width_adapter_003:in_ready -> id_router_003:src_ready
	wire          width_adapter_003_src_endofpacket;                                                                     // width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                                           // width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                                   // width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [106:0] width_adapter_003_src_data;                                                                            // width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	wire          width_adapter_003_src_ready;                                                                           // rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	wire   [10:0] width_adapter_003_src_channel;                                                                         // width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	wire          crosser_out_endofpacket;                                                                               // crosser:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                     // crosser:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                             // crosser:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] crosser_out_data;                                                                                      // crosser:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] crosser_out_channel;                                                                                   // crosser:out_channel -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                   // cmd_xbar_demux_001:src4_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                         // cmd_xbar_demux_001:src4_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                 // cmd_xbar_demux_001:src4_startofpacket -> crosser:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src4_data;                                                                          // cmd_xbar_demux_001:src4_data -> crosser:in_data
	wire   [10:0] cmd_xbar_demux_001_src4_channel;                                                                       // cmd_xbar_demux_001:src4_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                         // crosser:in_ready -> cmd_xbar_demux_001:src4_ready
	wire          crosser_001_out_endofpacket;                                                                           // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          crosser_001_out_valid;                                                                                 // crosser_001:out_valid -> rsp_xbar_mux_001:sink4_valid
	wire          crosser_001_out_startofpacket;                                                                         // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [106:0] crosser_001_out_data;                                                                                  // crosser_001:out_data -> rsp_xbar_mux_001:sink4_data
	wire   [10:0] crosser_001_out_channel;                                                                               // crosser_001:out_channel -> rsp_xbar_mux_001:sink4_channel
	wire          crosser_001_out_ready;                                                                                 // rsp_xbar_mux_001:sink4_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                   // rsp_xbar_demux_004:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                         // rsp_xbar_demux_004:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                 // rsp_xbar_demux_004:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                          // rsp_xbar_demux_004:src0_data -> crosser_001:in_data
	wire   [10:0] rsp_xbar_demux_004_src0_channel;                                                                       // rsp_xbar_demux_004:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                         // crosser_001:in_ready -> rsp_xbar_demux_004:src0_ready
	wire   [10:0] limiter_cmd_valid_data;                                                                                // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [10:0] limiter_001_cmd_valid_data;                                                                            // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire    [7:0] limiter_002_cmd_valid_data;                                                                            // limiter_002:cmd_src_valid -> cmd_xbar_demux_005:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                              // sgdma_pixel:csr_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                              // fifo:wrclk_control_slave_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                              // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                         // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver3_irq;                                                                              // irq_synchronizer:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                         // sys_clk_timer:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver4_irq;                                                                              // irq_synchronizer_001:sender_irq -> irq_mapper:receiver4_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                     // touch_panel_spi:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver5_irq;                                                                              // irq_synchronizer_002:sender_irq -> irq_mapper:receiver5_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                                     // touch_panel_pen_irq_n:irq -> irq_synchronizer_002:receiver_irq

	nios_simple_pll pll (
		.clk       (clk_ext),                                                //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                         // inclk_interface_reset.reset
		.read      (pll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (pll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (pll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (pll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (pll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (pll_c0_out),                                             //                    c0.clk
		.c1        (pll_c1_out),                                             //                    c1.clk
		.c2        (pll_c2_out),                                             //                    c2.clk
		.c3        (pll_c3_out),                                             //                    c3.clk
		.locked    (locked_from_the_pll),                                    //        locked_conduit.export
		.phasedone (phasedone_from_the_pll)                                  //     phasedone_conduit.export
	);

	nios_simple_sdram sdram (
		.clk            (pll_c2_out),                                            //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (zs_addr_from_the_sdram),                                //  wire.export
		.zs_ba          (zs_ba_from_the_sdram),                                  //      .export
		.zs_cas_n       (zs_cas_n_from_the_sdram),                               //      .export
		.zs_cke         (zs_cke_from_the_sdram),                                 //      .export
		.zs_cs_n        (zs_cs_n_from_the_sdram),                                //      .export
		.zs_dq          (zs_dq_to_and_from_the_sdram),                           //      .export
		.zs_dqm         (zs_dqm_from_the_sdram),                                 //      .export
		.zs_ras_n       (zs_ras_n_from_the_sdram),                               //      .export
		.zs_we_n        (zs_we_n_from_the_sdram)                                 //      .export
	);

	nios_simple_sgdma_pixel sgdma_pixel (
		.clk                           (pll_c2_out),                                                //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),                       //            reset.reset_n
		.csr_chipselect                (sgdma_pixel_csr_translator_avalon_anti_slave_0_chipselect), //              csr.chipselect
		.csr_address                   (sgdma_pixel_csr_translator_avalon_anti_slave_0_address),    //                 .address
		.csr_read                      (sgdma_pixel_csr_translator_avalon_anti_slave_0_read),       //                 .read
		.csr_write                     (sgdma_pixel_csr_translator_avalon_anti_slave_0_write),      //                 .write
		.csr_writedata                 (sgdma_pixel_csr_translator_avalon_anti_slave_0_writedata),  //                 .writedata
		.csr_readdata                  (sgdma_pixel_csr_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_pixel_descriptor_read_readdata),                      //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_pixel_descriptor_read_readdatavalid),                 //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_pixel_descriptor_read_waitrequest),                   //                 .waitrequest
		.descriptor_read_address       (sgdma_pixel_descriptor_read_address),                       //                 .address
		.descriptor_read_read          (sgdma_pixel_descriptor_read_read),                          //                 .read
		.descriptor_write_waitrequest  (sgdma_pixel_descriptor_write_waitrequest),                  // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_pixel_descriptor_write_address),                      //                 .address
		.descriptor_write_write        (sgdma_pixel_descriptor_write_write),                        //                 .write
		.descriptor_write_writedata    (sgdma_pixel_descriptor_write_writedata),                    //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                                  //          csr_irq.irq
		.m_read_readdata               (sgdma_pixel_m_read_readdata),                               //           m_read.readdata
		.m_read_readdatavalid          (sgdma_pixel_m_read_readdatavalid),                          //                 .readdatavalid
		.m_read_waitrequest            (sgdma_pixel_m_read_waitrequest),                            //                 .waitrequest
		.m_read_address                (sgdma_pixel_m_read_address),                                //                 .address
		.m_read_read                   (sgdma_pixel_m_read_read),                                   //                 .read
		.out_data                      (sgdma_pixel_out_data),                                      //              out.data
		.out_valid                     (sgdma_pixel_out_valid),                                     //                 .valid
		.out_ready                     (sgdma_pixel_out_ready),                                     //                 .ready
		.out_endofpacket               (sgdma_pixel_out_endofpacket),                               //                 .endofpacket
		.out_startofpacket             (sgdma_pixel_out_startofpacket),                             //                 .startofpacket
		.out_empty                     (sgdma_pixel_out_empty)                                      //                 .empty
	);

	nios_simple_fifo fifo (
		.wrclock                       (pll_c2_out),                                           //    clk_in.clk
		.wrreset_n                     (~rst_controller_001_reset_out_reset),                  //  reset_in.reset_n
		.rdclock                       (pll_c1_out),                                           //   clk_out.clk
		.rdreset_n                     (~rst_controller_002_reset_out_reset),                  // reset_out.reset_n
		.avalonst_sink_valid           (timing_adapter_out_valid),                             //        in.valid
		.avalonst_sink_data            (timing_adapter_out_data),                              //          .data
		.avalonst_sink_startofpacket   (timing_adapter_out_startofpacket),                     //          .startofpacket
		.avalonst_sink_endofpacket     (timing_adapter_out_endofpacket),                       //          .endofpacket
		.avalonst_sink_empty           (timing_adapter_out_empty),                             //          .empty
		.avalonst_sink_ready           (timing_adapter_out_ready),                             //          .ready
		.avalonst_source_valid         (fifo_out_valid),                                       //       out.valid
		.avalonst_source_data          (fifo_out_data),                                        //          .data
		.avalonst_source_startofpacket (fifo_out_startofpacket),                               //          .startofpacket
		.avalonst_source_endofpacket   (fifo_out_endofpacket),                                 //          .endofpacket
		.avalonst_source_empty         (fifo_out_empty),                                       //          .empty
		.avalonst_source_ready         (fifo_out_ready),                                       //          .ready
		.wrclk_control_slave_address   (fifo_in_csr_translator_avalon_anti_slave_0_address),   //    in_csr.address
		.wrclk_control_slave_read      (fifo_in_csr_translator_avalon_anti_slave_0_read),      //          .read
		.wrclk_control_slave_writedata (fifo_in_csr_translator_avalon_anti_slave_0_writedata), //          .writedata
		.wrclk_control_slave_write     (fifo_in_csr_translator_avalon_anti_slave_0_write),     //          .write
		.wrclk_control_slave_readdata  (fifo_in_csr_translator_avalon_anti_slave_0_readdata),  //          .readdata
		.wrclk_control_slave_irq       (irq_mapper_receiver1_irq)                              //    in_irq.irq
	);

	nios_simple_timing_adapter timing_adapter (
		.clk               (pll_c2_out),                          //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset), // reset.reset_n
		.in_ready          (sgdma_pixel_out_ready),               //    in.ready
		.in_valid          (sgdma_pixel_out_valid),               //      .valid
		.in_data           (sgdma_pixel_out_data),                //      .data
		.in_startofpacket  (sgdma_pixel_out_startofpacket),       //      .startofpacket
		.in_endofpacket    (sgdma_pixel_out_endofpacket),         //      .endofpacket
		.in_empty          (sgdma_pixel_out_empty),               //      .empty
		.out_ready         (timing_adapter_out_ready),            //   out.ready
		.out_valid         (timing_adapter_out_valid),            //      .valid
		.out_data          (timing_adapter_out_data),             //      .data
		.out_startofpacket (timing_adapter_out_startofpacket),    //      .startofpacket
		.out_endofpacket   (timing_adapter_out_endofpacket),      //      .endofpacket
		.out_empty         (timing_adapter_out_empty)             //      .empty
	);

	altera_avalon_pixel_converter pixel_converter (
		.clk       (pll_c1_out),                                //       clk.clk
		.reset_n   (~rst_controller_002_reset_out_reset),       // clk_reset.reset_n
		.ready_out (fifo_to_pixel_converter_out_ready),         //        in.ready
		.valid_in  (fifo_to_pixel_converter_out_valid),         //          .valid
		.data_in   (fifo_to_pixel_converter_out_data),          //          .data
		.eop_in    (fifo_to_pixel_converter_out_endofpacket),   //          .endofpacket
		.sop_in    (fifo_to_pixel_converter_out_startofpacket), //          .startofpacket
		.empty_in  (fifo_to_pixel_converter_out_empty),         //          .empty
		.ready_in  (pixel_converter_out_ready),                 //       out.ready
		.valid_out (pixel_converter_out_valid),                 //          .valid
		.data_out  (pixel_converter_out_data),                  //          .data
		.eop_out   (pixel_converter_out_endofpacket),           //          .endofpacket
		.sop_out   (pixel_converter_out_startofpacket),         //          .startofpacket
		.empty_out (pixel_converter_out_empty)                  //          .empty
	);

	altera_avalon_video_sync_generator video_sync_generator (
		.clk     (pll_c1_out),                            //       clk.clk
		.reset_n (~rst_controller_002_reset_out_reset),   // clk_reset.reset_n
		.ready   (pixel_converter_out_ready),             //        in.ready
		.valid   (pixel_converter_out_valid),             //          .valid
		.data    (pixel_converter_out_data),              //          .data
		.eop     (pixel_converter_out_endofpacket),       //          .endofpacket
		.sop     (pixel_converter_out_startofpacket),     //          .startofpacket
		.empty   (pixel_converter_out_empty),             //          .empty
		.RGB_OUT (RGB_OUT_from_the_video_sync_generator), //      sync.export
		.HD      (HD_from_the_video_sync_generator),      //          .export
		.VD      (VD_from_the_video_sync_generator),      //          .export
		.DEN     (DEN_from_the_video_sync_generator)      //          .export
	);

	nios_simple_fifo_to_pixel_converter fifo_to_pixel_converter (
		.clk               (pll_c1_out),                                //   clk.clk
		.reset_n           (~rst_controller_002_reset_out_reset),       // reset.reset_n
		.in_ready          (fifo_out_ready),                            //    in.ready
		.in_valid          (fifo_out_valid),                            //      .valid
		.in_data           (fifo_out_data),                             //      .data
		.in_startofpacket  (fifo_out_startofpacket),                    //      .startofpacket
		.in_endofpacket    (fifo_out_endofpacket),                      //      .endofpacket
		.in_empty          (fifo_out_empty),                            //      .empty
		.out_ready         (fifo_to_pixel_converter_out_ready),         //   out.ready
		.out_valid         (fifo_to_pixel_converter_out_valid),         //      .valid
		.out_data          (fifo_to_pixel_converter_out_data),          //      .data
		.out_startofpacket (fifo_to_pixel_converter_out_startofpacket), //      .startofpacket
		.out_endofpacket   (fifo_to_pixel_converter_out_endofpacket),   //      .endofpacket
		.out_empty         (fifo_to_pixel_converter_out_empty)          //      .empty
	);

	nios_simple_jtag_uart jtag_uart (
		.clk            (pll_c2_out),                                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                                //               irq.irq
	);

	sd_controller #(
		.IDLE                 (0),
		.SHIFT_OUT_CMD        (1),
		.WAIT_FOR_RSP_START   (2),
		.SHIFT_IN_CMD_RSP     (3),
		.WAIT_FOR_DATA_START  (4),
		.SHIFT_IN_DATA        (5),
		.SHIFT_IN_CRC16       (6),
		.SHIFT_OUT_DATA_TOKEN (7),
		.SHIFT_OUT_DATA       (8),
		.SHIFT_OUT_CRC16      (9),
		.SHIFT_IN_DATA_RSP    (10),
		.DATA_BUSY            (11),
		.ERROR_STATE          (12),
		.WAIT                 (13)
	) sd_card_controller (
		.clk                     (pll_c3_out),                                                                //       global_signals_clock.clk
		.reset_n                 (~rst_controller_003_reset_out_reset),                                       // global_signals_clock_reset.reset_n
		.avalon_slave_address    (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_address),    //               avalon_slave.address
		.avalon_slave_readdata   (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_readdata),   //                           .readdata
		.avalon_slave_writedata  (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_writedata),  //                           .writedata
		.avalon_slave_write      (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_write),      //                           .write
		.avalon_slave_read       (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_read),       //                           .read
		.avalon_slave_chipselect (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_chipselect), //                           .chipselect
		.avalon_slave_byteenable (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_byteenable), //                           .byteenable
		.spi_data_out            (spi_data_out_from_the_sd_card_controller),                                  //        avalon_slave_export.export
		.spi_data_in             (spi_data_in_to_the_sd_card_controller),                                     //                           .export
		.spi_cs_n                (spi_cs_n_from_the_sd_card_controller),                                      //                           .export
		.spi_clk                 (spi_clk_from_the_sd_card_controller)                                        //                           .export
	);

	nios_simple_lcd_i2c_scl lcd_i2c_scl (
		.clk        (pll_c3_out),                                               //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                      //               reset.reset_n
		.address    (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_i2c_scl_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_lcd_i2c_scl)                             // external_connection.export
	);

	nios_simple_lcd_i2c_scl lcd_i2c_en (
		.clk        (pll_c3_out),                                              //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                     //               reset.reset_n
		.address    (lcd_i2c_en_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_i2c_en_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_i2c_en_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_i2c_en_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_i2c_en_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (out_port_from_the_lcd_i2c_en)                             // external_connection.export
	);

	nios_simple_lcd_i2c_sda lcd_i2c_sda (
		.clk        (pll_c3_out),                                               //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                      //               reset.reset_n
		.address    (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~lcd_i2c_sda_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.bidir_port (bidir_port_to_and_from_the_lcd_i2c_sda)                    // external_connection.export
	);

	nios_simple_sys_clk_timer sys_clk_timer (
		.clk        (pll_c3_out),                                                 //   clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                        // reset.reset_n
		.address    (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_clk_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                               //   irq.irq
	);

	nios_simple_touch_panel_spi touch_panel_spi (
		.clk           (pll_c3_out),                                                                 //              clk.clk
		.reset_n       (~rst_controller_003_reset_out_reset),                                        //            reset.reset_n
		.data_from_cpu (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_writedata),  // spi_control_port.writedata
		.data_to_cpu   (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_readdata),   //                 .readdata
		.mem_addr      (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_address),    //                 .address
		.read_n        (~touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_read),      //                 .read_n
		.spi_select    (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_chipselect), //                 .chipselect
		.write_n       (~touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_write),     //                 .write_n
		.irq           (irq_synchronizer_001_receiver_irq),                                          //              irq.irq
		.MISO          (MISO_to_the_touch_panel_spi),                                                //         external.export
		.MOSI          (MOSI_from_the_touch_panel_spi),                                              //                 .export
		.SCLK          (SCLK_from_the_touch_panel_spi),                                              //                 .export
		.SS_n          (SS_n_from_the_touch_panel_spi)                                               //                 .export
	);

	nios_simple_touch_panel_pen_irq_n touch_panel_pen_irq_n (
		.clk        (pll_c3_out),                                                         //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),                                //               reset.reset_n
		.address    (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (in_port_to_the_touch_panel_pen_irq_n),                               // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)                                   //                 irq.irq
	);

	nios_simple_touch_panel_busy touch_panel_busy (
		.clk      (pll_c3_out),                                                  //                 clk.clk
		.reset_n  (~rst_controller_003_reset_out_reset),                         //               reset.reset_n
		.address  (touch_panel_busy_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (touch_panel_busy_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (in_port_to_the_touch_panel_busy)                              // external_connection.export
	);

	nios_simple_descriptor_mem descriptor_mem (
		.clk        (pll_c2_out),                                                  //   clk1.clk
		.address    (descriptor_mem_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (descriptor_mem_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (descriptor_mem_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (descriptor_mem_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (descriptor_mem_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (descriptor_mem_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (descriptor_mem_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                          // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)                       //       .reset_req
	);

	TERASIC_SRAM #(
		.DATA_BITS (16),
		.ADDR_BITS (20)
	) sram (
		.clk            (pll_c2_out),                                                   //       clock_reset.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                          // clock_reset_reset.reset_n
		.s_chipselect_n (~sram_avalon_slave_translator_avalon_anti_slave_0_chipselect), //      avalon_slave.chipselect_n
		.s_write_n      (~sram_avalon_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.s_address      (sram_avalon_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.s_read_n       (~sram_avalon_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.s_writedata    (sram_avalon_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.s_readdata     (sram_avalon_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.s_byteenable_n (~sram_avalon_slave_translator_avalon_anti_slave_0_byteenable), //                  .byteenable_n
		.SRAM_DQ        (SRAM_DQ_to_and_from_the_sram),                                 //       conduit_end.export
		.SRAM_ADDR      (SRAM_ADDR_from_the_sram),                                      //                  .export
		.SRAM_UB_n      (SRAM_UB_n_from_the_sram),                                      //                  .export
		.SRAM_LB_n      (SRAM_LB_n_from_the_sram),                                      //                  .export
		.SRAM_WE_n      (SRAM_WE_n_from_the_sram),                                      //                  .export
		.SRAM_CE_n      (SRAM_CE_n_from_the_sram),                                      //                  .export
		.SRAM_OE_n      (SRAM_OE_n_from_the_sram)                                       //                  .export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (11),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) peripheral_bridge (
		.m0_clk           (pll_c3_out),                                                        //   m0_clk.clk
		.m0_reset         (rst_controller_003_reset_out_reset),                                // m0_reset.reset
		.s0_clk           (pll_c2_out),                                                        //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                                // s0_reset.reset
		.s0_waitrequest   (peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (peripheral_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (peripheral_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (peripheral_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (peripheral_bridge_m0_address),                                      //         .address
		.m0_write         (peripheral_bridge_m0_write),                                        //         .write
		.m0_read          (peripheral_bridge_m0_read),                                         //         .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	nios_simple_cpu cpu (
		.clk                                   (pll_c2_out),                                                       //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                              //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                  // custom_instruction_master.readra
	);

	nios_simple_sysid sysid (
		.clock    (pll_c2_out),                                                  //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	nios_simple_tri_state_bridge_flash_bridge_0 tri_state_bridge_flash_bridge_0 (
		.clk                                   (pll_c2_out),                                                                //   clk.clk
		.reset                                 (rst_controller_001_reset_out_reset),                                        // reset.reset
		.request                               (tri_state_bridge_flash_pinsharer_0_tcm_request),                            //   tcs.request
		.grant                                 (tri_state_bridge_flash_pinsharer_0_tcm_grant),                              //      .grant
		.tcs_tri_state_bridge_flash_data       (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_out),    //      .tri_state_bridge_flash_data_out
		.tcs_tri_state_bridge_flash_data_outen (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_outen),  //      .tri_state_bridge_flash_data_outen
		.tcs_tri_state_bridge_flash_data_in    (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_in),     //      .tri_state_bridge_flash_data_in
		.tcs_write_n_to_the_cfi_flash          (tri_state_bridge_flash_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),       //      .write_n_to_the_cfi_flash_out
		.tcs_select_n_to_the_cfi_flash         (tri_state_bridge_flash_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),      //      .select_n_to_the_cfi_flash_out
		.tcs_read_n_to_the_cfi_flash           (tri_state_bridge_flash_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),        //      .read_n_to_the_cfi_flash_out
		.tcs_tri_state_bridge_flash_address    (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_address_out), //      .tri_state_bridge_flash_address_out
		.tri_state_bridge_flash_data           (tri_state_bridge_flash_data),                                               //   out.tri_state_bridge_flash_data
		.write_n_to_the_cfi_flash              (write_n_to_the_cfi_flash),                                                  //      .write_n_to_the_cfi_flash
		.select_n_to_the_cfi_flash             (select_n_to_the_cfi_flash),                                                 //      .select_n_to_the_cfi_flash
		.read_n_to_the_cfi_flash               (read_n_to_the_cfi_flash),                                                   //      .read_n_to_the_cfi_flash
		.tri_state_bridge_flash_address        (tri_state_bridge_flash_address)                                             //      .tri_state_bridge_flash_address
	);

	nios_simple_tri_state_bridge_flash_pinSharer_0 tri_state_bridge_flash_pinsharer_0 (
		.clk_clk                           (pll_c2_out),                                                                //   clk.clk
		.reset_reset                       (rst_controller_001_reset_out_reset),                                        // reset.reset
		.request                           (tri_state_bridge_flash_pinsharer_0_tcm_request),                            //   tcm.request
		.grant                             (tri_state_bridge_flash_pinsharer_0_tcm_grant),                              //      .grant
		.tri_state_bridge_flash_address    (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_address_out), //      .tri_state_bridge_flash_address_out
		.read_n_to_the_cfi_flash           (tri_state_bridge_flash_pinsharer_0_tcm_read_n_to_the_cfi_flash_out),        //      .read_n_to_the_cfi_flash_out
		.write_n_to_the_cfi_flash          (tri_state_bridge_flash_pinsharer_0_tcm_write_n_to_the_cfi_flash_out),       //      .write_n_to_the_cfi_flash_out
		.tri_state_bridge_flash_data       (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_out),    //      .tri_state_bridge_flash_data_out
		.tri_state_bridge_flash_data_in    (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_in),     //      .tri_state_bridge_flash_data_in
		.tri_state_bridge_flash_data_outen (tri_state_bridge_flash_pinsharer_0_tcm_tri_state_bridge_flash_data_outen),  //      .tri_state_bridge_flash_data_outen
		.select_n_to_the_cfi_flash         (tri_state_bridge_flash_pinsharer_0_tcm_select_n_to_the_cfi_flash_out),      //      .select_n_to_the_cfi_flash_out
		.tcs0_request                      (cfi_flash_tcm_request),                                                     //  tcs0.request
		.tcs0_grant                        (cfi_flash_tcm_grant),                                                       //      .grant
		.tcs0_address_out                  (cfi_flash_tcm_address_out),                                                 //      .address_out
		.tcs0_read_n_out                   (cfi_flash_tcm_read_n_out),                                                  //      .read_n_out
		.tcs0_write_n_out                  (cfi_flash_tcm_write_n_out),                                                 //      .write_n_out
		.tcs0_data_out                     (cfi_flash_tcm_data_out),                                                    //      .data_out
		.tcs0_data_in                      (cfi_flash_tcm_data_in),                                                     //      .data_in
		.tcs0_data_outen                   (cfi_flash_tcm_data_outen),                                                  //      .data_outen
		.tcs0_chipselect_n_out             (cfi_flash_tcm_chipselect_n_out)                                             //      .chipselect_n_out
	);

	nios_simple_cfi_flash #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (60),
		.TCM_DATA_HOLD                  (60),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) cfi_flash (
		.clk_clk              (pll_c2_out),                                                 //   clk.clk
		.reset_reset          (rst_controller_001_reset_out_reset),                         // reset.reset
		.uas_address          (cfi_flash_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (cfi_flash_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (cfi_flash_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (cfi_flash_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (cfi_flash_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (cfi_flash_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (cfi_flash_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (cfi_flash_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (cfi_flash_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (cfi_flash_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (cfi_flash_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (cfi_flash_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (cfi_flash_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (cfi_flash_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (cfi_flash_tcm_request),                                      //      .request
		.tcm_grant            (cfi_flash_tcm_grant),                                        //      .grant
		.tcm_address_out      (cfi_flash_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (cfi_flash_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (cfi_flash_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (cfi_flash_tcm_data_in)                                       //      .data_in
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                      (pll_c2_out),                                                                //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                        //                     reset.reset
		.uav_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_byteenable            (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_write                 (1'b0),                                                                      //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (28),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                      (pll_c2_out),                                                         //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address              (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_data_master_read),                                               //                          .read
		.av_readdata              (cpu_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (cpu_data_master_write),                                              //                          .write
		.av_writedata             (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_pixel_descriptor_write_translator (
		.clk                      (pll_c2_out),                                                                      //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                              //                     reset.reset
		.uav_address              (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (sgdma_pixel_descriptor_write_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (sgdma_pixel_descriptor_write_waitrequest),                                        //                          .waitrequest
		.av_write                 (sgdma_pixel_descriptor_write_write),                                              //                          .write
		.av_writedata             (sgdma_pixel_descriptor_write_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                            //               (terminated)
		.av_byteenable            (4'b1111),                                                                         //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                            //               (terminated)
		.av_begintransfer         (1'b0),                                                                            //               (terminated)
		.av_chipselect            (1'b0),                                                                            //               (terminated)
		.av_read                  (1'b0),                                                                            //               (terminated)
		.av_readdata              (),                                                                                //               (terminated)
		.av_readdatavalid         (),                                                                                //               (terminated)
		.av_lock                  (1'b0),                                                                            //               (terminated)
		.av_debugaccess           (1'b0),                                                                            //               (terminated)
		.uav_clken                (),                                                                                //               (terminated)
		.av_clken                 (1'b1),                                                                            //               (terminated)
		.uav_response             (2'b00),                                                                           //               (terminated)
		.av_response              (),                                                                                //               (terminated)
		.uav_writeresponserequest (),                                                                                //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                            //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                            //               (terminated)
		.av_writeresponsevalid    ()                                                                                 //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_pixel_descriptor_read_translator (
		.clk                      (pll_c2_out),                                                                     //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                     reset.reset
		.uav_address              (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (sgdma_pixel_descriptor_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (sgdma_pixel_descriptor_read_waitrequest),                                        //                          .waitrequest
		.av_read                  (sgdma_pixel_descriptor_read_read),                                               //                          .read
		.av_readdata              (sgdma_pixel_descriptor_read_readdata),                                           //                          .readdata
		.av_readdatavalid         (sgdma_pixel_descriptor_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                           //               (terminated)
		.av_byteenable            (4'b1111),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                           //               (terminated)
		.av_begintransfer         (1'b0),                                                                           //               (terminated)
		.av_chipselect            (1'b0),                                                                           //               (terminated)
		.av_write                 (1'b0),                                                                           //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                           //               (terminated)
		.av_lock                  (1'b0),                                                                           //               (terminated)
		.av_debugaccess           (1'b0),                                                                           //               (terminated)
		.uav_clken                (),                                                                               //               (terminated)
		.av_clken                 (1'b1),                                                                           //               (terminated)
		.uav_response             (2'b00),                                                                          //               (terminated)
		.av_response              (),                                                                               //               (terminated)
		.uav_writeresponserequest (),                                                                               //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                           //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                           //               (terminated)
		.av_writeresponsevalid    ()                                                                                //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) sgdma_pixel_m_read_translator (
		.clk                      (pll_c2_out),                                                            //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                     reset.reset
		.uav_address              (sgdma_pixel_m_read_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (sgdma_pixel_m_read_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (sgdma_pixel_m_read_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (sgdma_pixel_m_read_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (sgdma_pixel_m_read_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (sgdma_pixel_m_read_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (sgdma_pixel_m_read_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (sgdma_pixel_m_read_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (sgdma_pixel_m_read_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (sgdma_pixel_m_read_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (sgdma_pixel_m_read_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (sgdma_pixel_m_read_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (sgdma_pixel_m_read_waitrequest),                                        //                          .waitrequest
		.av_read                  (sgdma_pixel_m_read_read),                                               //                          .read
		.av_readdata              (sgdma_pixel_m_read_readdata),                                           //                          .readdata
		.av_readdatavalid         (sgdma_pixel_m_read_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                  //               (terminated)
		.av_byteenable            (4'b1111),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                  //               (terminated)
		.av_chipselect            (1'b0),                                                                  //               (terminated)
		.av_write                 (1'b0),                                                                  //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                  //               (terminated)
		.av_lock                  (1'b0),                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                  //               (terminated)
		.uav_clken                (),                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                 //               (terminated)
		.av_response              (),                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                      (pll_c2_out),                                                                       //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                               //                    reset.reset
		.uav_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (2),
		.AV_SETUP_WAIT_CYCLES           (1),
		.AV_DATA_HOLD_CYCLES            (1)
	) sram_avalon_slave_translator (
		.clk                      (pll_c2_out),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sram_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sram_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sram_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sram_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sram_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sram_avalon_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (sram_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (pll_c2_out),                                                          //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (23),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cfi_flash_uas_translator (
		.clk                      (pll_c2_out),                                                               //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                       //                    reset.reset
		.uav_address              (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cfi_flash_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cfi_flash_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cfi_flash_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cfi_flash_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cfi_flash_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (cfi_flash_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (cfi_flash_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (cfi_flash_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (cfi_flash_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock                  (cfi_flash_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess           (cfi_flash_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_chipselect            (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pll_pll_slave_translator (
		.clk                      (clk_ext),                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_chipselect            (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sgdma_pixel_csr_translator (
		.clk                      (pll_c2_out),                                                                 //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                         //                    reset.reset
		.uav_address              (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sgdma_pixel_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sgdma_pixel_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sgdma_pixel_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sgdma_pixel_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sgdma_pixel_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sgdma_pixel_csr_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_byteenable            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fifo_in_csr_translator (
		.clk                      (pll_c2_out),                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                     //                    reset.reset
		.uav_address              (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fifo_in_csr_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fifo_in_csr_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fifo_in_csr_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fifo_in_csr_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fifo_in_csr_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (pll_c2_out),                                                                             //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (pll_c2_out),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (14),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) descriptor_mem_s1_translator (
		.clk                      (pll_c2_out),                                                                   //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                           //                    reset.reset
		.uav_address              (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (descriptor_mem_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (descriptor_mem_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (descriptor_mem_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (descriptor_mem_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (descriptor_mem_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (descriptor_mem_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (descriptor_mem_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) peripheral_bridge_s0_translator (
		.clk                      (pll_c2_out),                                                                      //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                              //                    reset.reset
		.uav_address              (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (peripheral_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (peripheral_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (peripheral_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.av_chipselect            (),                                                                                //              (terminated)
		.av_clken                 (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (11),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (11),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) peripheral_bridge_m0_translator (
		.clk                      (pll_c3_out),                                                              //                       clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                      //                     reset.reset
		.uav_address              (peripheral_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (peripheral_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (peripheral_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (peripheral_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (peripheral_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (peripheral_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (peripheral_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (peripheral_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (peripheral_bridge_m0_read),                                               //                          .read
		.av_readdata              (peripheral_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (peripheral_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (peripheral_bridge_m0_write),                                              //                          .write
		.av_writedata             (peripheral_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (peripheral_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                    //               (terminated)
		.av_lock                  (1'b0),                                                                    //               (terminated)
		.uav_clken                (),                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                   //               (terminated)
		.av_response              (),                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sd_card_controller_avalon_slave_translator (
		.clk                      (pll_c3_out),                                                                                 //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (sd_card_controller_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                                           //              (terminated)
		.av_burstcount            (),                                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                                           //              (terminated)
		.av_lock                  (),                                                                                           //              (terminated)
		.av_clken                 (),                                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                                       //              (terminated)
		.av_debugaccess           (),                                                                                           //              (terminated)
		.av_outputenable          (),                                                                                           //              (terminated)
		.uav_response             (),                                                                                           //              (terminated)
		.av_response              (2'b00),                                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_i2c_scl_s1_translator (
		.clk                      (pll_c3_out),                                                                //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                        //                    reset.reset
		.uav_address              (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_i2c_scl_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_i2c_en_s1_translator (
		.clk                      (pll_c3_out),                                                               //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                       //                    reset.reset
		.uav_address              (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_i2c_en_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_i2c_en_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_i2c_en_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_i2c_en_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_i2c_en_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) lcd_i2c_sda_s1_translator (
		.clk                      (pll_c3_out),                                                                //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                        //                    reset.reset
		.uav_address              (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (lcd_i2c_sda_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                          //              (terminated)
		.av_begintransfer         (),                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                          //              (terminated)
		.av_burstcount            (),                                                                          //              (terminated)
		.av_byteenable            (),                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                      //              (terminated)
		.av_waitrequest           (1'b0),                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                          //              (terminated)
		.av_lock                  (),                                                                          //              (terminated)
		.av_clken                 (),                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                      //              (terminated)
		.av_debugaccess           (),                                                                          //              (terminated)
		.av_outputenable          (),                                                                          //              (terminated)
		.uav_response             (),                                                                          //              (terminated)
		.av_response              (2'b00),                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_clk_timer_s1_translator (
		.clk                      (pll_c3_out),                                                                  //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                          //                    reset.reset
		.uav_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sys_clk_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) touch_panel_spi_spi_control_port_translator (
		.clk                      (pll_c3_out),                                                                                  //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (touch_panel_spi_spi_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                                            //              (terminated)
		.av_burstcount            (),                                                                                            //              (terminated)
		.av_byteenable            (),                                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                                            //              (terminated)
		.av_lock                  (),                                                                                            //              (terminated)
		.av_clken                 (),                                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                                        //              (terminated)
		.av_debugaccess           (),                                                                                            //              (terminated)
		.av_outputenable          (),                                                                                            //              (terminated)
		.uav_response             (),                                                                                            //              (terminated)
		.av_response              (2'b00),                                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) touch_panel_pen_irq_n_s1_translator (
		.clk                      (pll_c3_out),                                                                          //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (touch_panel_pen_irq_n_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                    //              (terminated)
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (11),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) touch_panel_busy_s1_translator (
		.clk                      (pll_c3_out),                                                                     //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                             //                    reset.reset
		.uav_address              (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (touch_panel_busy_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (touch_panel_busy_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c2_out),                                                                         //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.av_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                              //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                               //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                            //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                      //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                        //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                              //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c2_out),                                                                  //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address              (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                   //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                    //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                 //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                           //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                             //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                   //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c2_out),                                                                               //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_009_src1_valid),                                                            //        rp.valid
		.rp_data                 (rsp_xbar_demux_009_src1_data),                                                             //          .data
		.rp_channel              (rsp_xbar_demux_009_src1_channel),                                                          //          .channel
		.rp_startofpacket        (rsp_xbar_demux_009_src1_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_009_src1_endofpacket),                                                      //          .endofpacket
		.rp_ready                (rsp_xbar_demux_009_src1_ready),                                                            //          .ready
		.av_response             (),                                                                                         // (terminated)
		.av_writeresponserequest (1'b0),                                                                                     // (terminated)
		.av_writeresponsevalid   ()                                                                                          // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c2_out),                                                                              //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.av_address              (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_009_src2_valid),                                                           //        rp.valid
		.rp_data                 (rsp_xbar_demux_009_src2_data),                                                            //          .data
		.rp_channel              (rsp_xbar_demux_009_src2_channel),                                                         //          .channel
		.rp_startofpacket        (rsp_xbar_demux_009_src2_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_009_src2_endofpacket),                                                     //          .endofpacket
		.rp_ready                (rsp_xbar_demux_009_src2_ready),                                                           //          .ready
		.av_response             (),                                                                                        // (terminated)
		.av_writeresponserequest (1'b0),                                                                                    // (terminated)
		.av_writeresponsevalid   ()                                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_pixel_m_read_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c2_out),                                                                     //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.av_address              (sgdma_pixel_m_read_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (sgdma_pixel_m_read_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (sgdma_pixel_m_read_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (sgdma_pixel_m_read_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (sgdma_pixel_m_read_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (sgdma_pixel_m_read_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (sgdma_pixel_m_read_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (sgdma_pixel_m_read_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (sgdma_pixel_m_read_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (sgdma_pixel_m_read_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (sgdma_pixel_m_read_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_002_src2_valid),                                                  //        rp.valid
		.rp_data                 (rsp_xbar_demux_002_src2_data),                                                   //          .data
		.rp_channel              (rsp_xbar_demux_002_src2_channel),                                                //          .channel
		.rp_startofpacket        (rsp_xbar_demux_002_src2_startofpacket),                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_002_src2_endofpacket),                                            //          .endofpacket
		.rp_ready                (rsp_xbar_demux_002_src2_ready),                                                  //          .ready
		.av_response             (),                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                   //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sram_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sram_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                            //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                            //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                             //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                          //                .channel
		.rf_sink_ready           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                  //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (65),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (66),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cfi_flash_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cfi_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                    //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                    //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                     //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                  //                .channel
		.rf_sink_ready           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (10),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c2_out),                                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.in_data           (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_ext),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                  //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                  //                .valid
		.cp_data                 (crosser_out_data),                                                                   //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                            //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                //                .channel
		.rf_sink_ready           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_ext),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_ext),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sgdma_pixel_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                           //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                      //                .channel
		.rf_sink_ready           (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fifo_in_csr_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fifo_in_csr_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                  //                .channel
		.rf_sink_ready           (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fifo_in_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.in_data           (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fifo_in_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fifo_in_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                       //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                       //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) descriptor_mem_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                             //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                             //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                             //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                              //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                       //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                           //                .channel
		.rf_sink_ready           (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                             //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) peripheral_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                          //                .channel
		.rf_sink_ready           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (97),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_BEGIN_BURST           (64),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.PKT_BURST_TYPE_H          (61),
		.PKT_BURST_TYPE_L          (60),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_TRANS_EXCLUSIVE       (52),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (72),
		.PKT_THREAD_ID_L           (72),
		.PKT_CACHE_H               (79),
		.PKT_CACHE_L               (76),
		.PKT_DATA_SIDEBAND_H       (63),
		.PKT_DATA_SIDEBAND_L       (63),
		.PKT_QOS_H                 (65),
		.PKT_QOS_L                 (65),
		.PKT_ADDR_SIDEBAND_H       (62),
		.PKT_ADDR_SIDEBAND_L       (62),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (8),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) peripheral_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c3_out),                                                                       //       clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.av_address              (peripheral_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (peripheral_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (peripheral_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (peripheral_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_002_rsp_src_valid),                                                        //        rp.valid
		.rp_data                 (limiter_002_rsp_src_data),                                                         //          .data
		.rp_channel              (limiter_002_rsp_src_channel),                                                      //          .channel
		.rp_startofpacket        (limiter_002_rsp_src_startofpacket),                                                //          .startofpacket
		.rp_endofpacket          (limiter_002_rsp_src_endofpacket),                                                  //          .endofpacket
		.rp_ready                (limiter_002_rsp_src_ready),                                                        //          .ready
		.av_response             (),                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                                           //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src0_ready),                                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src0_valid),                                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_005_src0_data),                                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src0_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src0_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src0_channel),                                                                      //                .channel
		.rf_sink_ready           (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                                           //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                                 // (terminated)
		.csr_readdata      (),                                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                 // (terminated)
		.almost_full_data  (),                                                                                                     // (terminated)
		.almost_empty_data (),                                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                                 // (terminated)
		.out_empty         (),                                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                                 // (terminated)
		.out_error         (),                                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                                 // (terminated)
		.out_channel       ()                                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                          //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src1_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src1_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_005_src1_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src1_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src1_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src1_channel),                                                     //                .channel
		.rf_sink_ready           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                         //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src2_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src2_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_005_src2_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src2_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src2_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src2_channel),                                                    //                .channel
		.rf_sink_ready           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                         //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                          //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src3_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src3_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_005_src3_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src3_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src3_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src3_channel),                                                     //                .channel
		.rf_sink_ready           (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                            //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src4_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src4_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_005_src4_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src4_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src4_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src4_channel),                                                       //                .channel
		.rf_sink_ready           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                                            //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src5_ready),                                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src5_valid),                                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_005_src5_data),                                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src5_startofpacket),                                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src5_endofpacket),                                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src5_channel),                                                                       //                .channel
		.rf_sink_ready           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                                    //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src6_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src6_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_005_src6_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src6_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src6_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src6_channel),                                                               //                .channel
		.rf_sink_ready           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                                    //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (64),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (46),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (47),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.PKT_TRANS_READ            (50),
		.PKT_TRANS_LOCK            (51),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (66),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (56),
		.PKT_BURSTWRAP_L           (56),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (59),
		.PKT_BURST_SIZE_L          (57),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) touch_panel_busy_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c3_out),                                                                               //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_005_src7_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_005_src7_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_005_src7_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_005_src7_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_005_src7_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_005_src7_channel),                                                          //                .channel
		.rf_sink_ready           (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c3_out),                                                                               //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	nios_simple_addr_router addr_router (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                              //       src.ready
		.src_valid          (addr_router_src_valid),                                                              //          .valid
		.src_data           (addr_router_src_data),                                                               //          .data
		.src_channel        (addr_router_src_channel),                                                            //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios_simple_addr_router_001 addr_router_001 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                  //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                              //          .endofpacket
	);

	nios_simple_addr_router_002 addr_router_002 (
		.sink_ready         (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_pixel_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                                //          .valid
		.src_data           (addr_router_002_src_data),                                                                 //          .data
		.src_channel        (addr_router_002_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                           //          .endofpacket
	);

	nios_simple_addr_router_002 addr_router_003 (
		.sink_ready         (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_pixel_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                              //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                               //          .valid
		.src_data           (addr_router_003_src_data),                                                                //          .data
		.src_channel        (addr_router_003_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                          //          .endofpacket
	);

	nios_simple_addr_router_004 addr_router_004 (
		.sink_ready         (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_pixel_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                      //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                      //          .valid
		.src_data           (addr_router_004_src_data),                                                       //          .data
		.src_channel        (addr_router_004_src_channel),                                                    //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                 //          .endofpacket
	);

	nios_simple_id_router id_router (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                              //       src.ready
		.src_valid          (id_router_src_valid),                                                              //          .valid
		.src_data           (id_router_src_data),                                                               //          .data
		.src_channel        (id_router_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                         //          .endofpacket
	);

	nios_simple_id_router_001 id_router_001 (
		.sink_ready         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sram_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                      //       src.ready
		.src_valid          (id_router_001_src_valid),                                                      //          .valid
		.src_data           (id_router_001_src_data),                                                       //          .data
		.src_channel        (id_router_001_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                 //          .endofpacket
	);

	nios_simple_id_router_002 id_router_002 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                             //       src.ready
		.src_valid          (id_router_002_src_valid),                                             //          .valid
		.src_data           (id_router_002_src_data),                                              //          .data
		.src_channel        (id_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                        //          .endofpacket
	);

	nios_simple_id_router_003 id_router_003 (
		.sink_ready         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cfi_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                  //       src.ready
		.src_valid          (id_router_003_src_valid),                                                  //          .valid
		.src_data           (id_router_003_src_data),                                                   //          .data
		.src_channel        (id_router_003_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                             //          .endofpacket
	);

	nios_simple_id_router_004 id_router_004 (
		.sink_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_ext),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                  //       src.ready
		.src_valid          (id_router_004_src_valid),                                                  //          .valid
		.src_data           (id_router_004_src_data),                                                   //          .data
		.src_channel        (id_router_004_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                             //          .endofpacket
	);

	nios_simple_id_router_004 id_router_005 (
		.sink_ready         (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sgdma_pixel_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                 //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                    //       src.ready
		.src_valid          (id_router_005_src_valid),                                                    //          .valid
		.src_data           (id_router_005_src_data),                                                     //          .data
		.src_channel        (id_router_005_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                               //          .endofpacket
	);

	nios_simple_id_router_004 id_router_006 (
		.sink_ready         (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fifo_in_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                //       src.ready
		.src_valid          (id_router_006_src_valid),                                                //          .valid
		.src_data           (id_router_006_src_data),                                                 //          .data
		.src_channel        (id_router_006_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                           //          .endofpacket
	);

	nios_simple_id_router_004 id_router_007 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                             //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                                //       src.ready
		.src_valid          (id_router_007_src_valid),                                                                //          .valid
		.src_data           (id_router_007_src_data),                                                                 //          .data
		.src_channel        (id_router_007_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                           //          .endofpacket
	);

	nios_simple_id_router_004 id_router_008 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                        //       src.ready
		.src_valid          (id_router_008_src_valid),                                                        //          .valid
		.src_data           (id_router_008_src_data),                                                         //          .data
		.src_channel        (id_router_008_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                   //          .endofpacket
	);

	nios_simple_id_router_009 id_router_009 (
		.sink_ready         (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (descriptor_mem_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                      //       src.ready
		.src_valid          (id_router_009_src_valid),                                                      //          .valid
		.src_data           (id_router_009_src_data),                                                       //          .data
		.src_channel        (id_router_009_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                 //          .endofpacket
	);

	nios_simple_id_router_004 id_router_010 (
		.sink_ready         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                         //       src.ready
		.src_valid          (id_router_010_src_valid),                                                         //          .valid
		.src_data           (id_router_010_src_data),                                                          //          .data
		.src_channel        (id_router_010_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                    //          .endofpacket
	);

	nios_simple_addr_router_005 addr_router_005 (
		.sink_ready         (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                       //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                        //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                        //          .valid
		.src_data           (addr_router_005_src_data),                                                         //          .data
		.src_channel        (addr_router_005_src_channel),                                                      //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                   //          .endofpacket
	);

	nios_simple_id_router_011 id_router_011 (
		.sink_ready         (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sd_card_controller_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                                 //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                                    //       src.ready
		.src_valid          (id_router_011_src_valid),                                                                    //          .valid
		.src_data           (id_router_011_src_data),                                                                     //          .data
		.src_channel        (id_router_011_src_channel),                                                                  //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                            //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                               //          .endofpacket
	);

	nios_simple_id_router_011 id_router_012 (
		.sink_ready         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_i2c_scl_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                   //       src.ready
		.src_valid          (id_router_012_src_valid),                                                   //          .valid
		.src_data           (id_router_012_src_data),                                                    //          .data
		.src_channel        (id_router_012_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                              //          .endofpacket
	);

	nios_simple_id_router_011 id_router_013 (
		.sink_ready         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_i2c_en_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                               //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                  //       src.ready
		.src_valid          (id_router_013_src_valid),                                                  //          .valid
		.src_data           (id_router_013_src_data),                                                   //          .data
		.src_channel        (id_router_013_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                             //          .endofpacket
	);

	nios_simple_id_router_011 id_router_014 (
		.sink_ready         (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_i2c_sda_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                   //       src.ready
		.src_valid          (id_router_014_src_valid),                                                   //          .valid
		.src_data           (id_router_014_src_data),                                                    //          .data
		.src_channel        (id_router_014_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                              //          .endofpacket
	);

	nios_simple_id_router_011 id_router_015 (
		.sink_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                     //       src.ready
		.src_valid          (id_router_015_src_valid),                                                     //          .valid
		.src_data           (id_router_015_src_data),                                                      //          .data
		.src_channel        (id_router_015_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                //          .endofpacket
	);

	nios_simple_id_router_011 id_router_016 (
		.sink_ready         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (touch_panel_spi_spi_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                                  //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_016_src_valid),                                                                     //          .valid
		.src_data           (id_router_016_src_data),                                                                      //          .data
		.src_channel        (id_router_016_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                                //          .endofpacket
	);

	nios_simple_id_router_011 id_router_017 (
		.sink_ready         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (touch_panel_pen_irq_n_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                          //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                             //       src.ready
		.src_valid          (id_router_017_src_valid),                                                             //          .valid
		.src_data           (id_router_017_src_data),                                                              //          .data
		.src_channel        (id_router_017_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                        //          .endofpacket
	);

	nios_simple_id_router_011 id_router_018 (
		.sink_ready         (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (touch_panel_busy_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c3_out),                                                                     //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                                        //       src.ready
		.src_valid          (id_router_018_src_valid),                                                        //          .valid
		.src_data           (id_router_018_src_data),                                                         //          .data
		.src_channel        (id_router_018_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                                   //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (11),
		.VALID_WIDTH               (11),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (pll_c2_out),                         //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),              //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),              //          .valid
		.cmd_sink_data          (addr_router_src_data),               //          .data
		.cmd_sink_channel       (addr_router_src_channel),            //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),             //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),             //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),           //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),              //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),     //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),       //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (96),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (11),
		.VALID_WIDTH               (11),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (pll_c2_out),                         //       clk.clk
		.reset                  (rst_controller_001_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (69),
		.PKT_TRANS_POSTED          (48),
		.PKT_TRANS_WRITE           (49),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (8),
		.VALID_WIDTH               (8),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (55),
		.PKT_BYTE_CNT_L            (53),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (pll_c3_out),                         //       clk.clk
		.reset                  (rst_controller_003_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_005_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_005_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_005_src_data),           //          .data
		.cmd_sink_channel       (addr_router_005_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_005_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_005_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_005_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_005_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_005_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_005_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_005_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_005_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (pll_c2_out),                          //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (11),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (pll_c2_out),                              //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_n),                          // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_ext),                           //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_req  (),                                  // (terminated)
		.reset_in2  (1'b0),                              // (terminated)
		.reset_in3  (1'b0),                              // (terminated)
		.reset_in4  (1'b0),                              // (terminated)
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller_001 (
		.reset_in0  (~reset_n),                               // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk        (pll_c2_out),                             //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_in2  (1'b0),                                   // (terminated)
		.reset_in3  (1'b0),                                   // (terminated)
		.reset_in4  (1'b0),                                   // (terminated)
		.reset_in5  (1'b0),                                   // (terminated)
		.reset_in6  (1'b0),                                   // (terminated)
		.reset_in7  (1'b0),                                   // (terminated)
		.reset_in8  (1'b0),                                   // (terminated)
		.reset_in9  (1'b0),                                   // (terminated)
		.reset_in10 (1'b0),                                   // (terminated)
		.reset_in11 (1'b0),                                   // (terminated)
		.reset_in12 (1'b0),                                   // (terminated)
		.reset_in13 (1'b0),                                   // (terminated)
		.reset_in14 (1'b0),                                   // (terminated)
		.reset_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (pll_c1_out),                         //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_003 (
		.reset_in0  (~reset_n),                           // reset_in0.reset
		.reset_in1  (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk        (pll_c3_out),                         //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_simple_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pll_c2_out),                         //        clk.clk
		.reset              (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),            //           .channel
		.sink_data          (limiter_cmd_src_data),               //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)     //           .endofpacket
	);

	nios_simple_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (pll_c2_out),                             //        clk.clk
		.reset               (rst_controller_001_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket)    //           .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 cmd_xbar_demux_003 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 cmd_xbar_demux_004 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (pll_c2_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (pll_c2_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (pll_c2_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (pll_c2_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_mux_009 cmd_xbar_mux_009 (
		.clk                 (pll_c2_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src9_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src9_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_003_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pll_c2_out),                         //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (id_router_src_ready),                //      sink.ready
		.sink_channel       (id_router_src_channel),              //          .channel
		.sink_data          (id_router_src_data),                 //          .data
		.sink_startofpacket (id_router_src_startofpacket),        //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),          //          .endofpacket
		.sink_valid         (id_router_src_valid),                //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),          //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),           //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),    //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),          //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),          //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),           //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),        //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)     //          .endofpacket
	);

	nios_simple_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_002_src2_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_ext),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_009_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_009_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_009_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_009_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_009_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_009_src2_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pll_c2_out),                            //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (pll_c2_out),                            //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (crosser_001_out_ready),                 //     sink4.ready
		.sink4_valid          (crosser_001_out_valid),                 //          .valid
		.sink4_channel        (crosser_001_out_channel),               //          .channel
		.sink4_data           (crosser_001_out_data),                  //          .data
		.sink4_startofpacket  (crosser_001_out_startofpacket),         //          .startofpacket
		.sink4_endofpacket    (crosser_001_out_endofpacket),           //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_cmd_xbar_demux_005 cmd_xbar_demux_005 (
		.clk                (pll_c3_out),                            //        clk.clk
		.reset              (rst_controller_003_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_005_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_005_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_005_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_005_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_005_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_005_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_005_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_005_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_005_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_005_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_005_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_005_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_005_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_005_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_005_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_005_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_005_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_005_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_005_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_005_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_005_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_005_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_005_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_005_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_005_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_005_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_005_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_005_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_005_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_005_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_005_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_005_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_005_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_005_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_005_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_005_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_005_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_005_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_005_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_005_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_005_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_005_src7_endofpacket)    //           .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_011 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_012 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_013 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_014 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_015 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_016 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_017 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_demux_011 rsp_xbar_demux_018 (
		.clk                (pll_c3_out),                            //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_simple_rsp_xbar_mux_005 rsp_xbar_mux_005 (
		.clk                 (pll_c3_out),                            //       clk.clk
		.reset               (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_005_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_005_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_011_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_012_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_013_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_014_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_015_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_016_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink6_ready         (rsp_xbar_demux_017_src0_ready),         //     sink6.ready
		.sink6_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink6_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink6_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink6_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink7_ready         (rsp_xbar_demux_018_src0_ready),         //     sink7.ready
		.sink7_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink7_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink7_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink7_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (pll_c2_out),                         //       clk.clk
		.reset                (rst_controller_001_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (pll_c2_out),                          //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (pll_c2_out),                          //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (cmd_xbar_mux_003_src_valid),          //      sink.valid
		.in_channel           (cmd_xbar_mux_003_src_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_mux_003_src_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_003_src_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_mux_003_src_ready),          //          .ready
		.in_data              (cmd_xbar_mux_003_src_data),           //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (11),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_003 (
		.clk                  (pll_c2_out),                          //       clk.clk
		.reset                (rst_controller_001_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_003_src_valid),             //      sink.valid
		.in_channel           (id_router_003_src_channel),           //          .channel
		.in_startofpacket     (id_router_003_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_003_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_003_src_ready),             //          .ready
		.in_data              (id_router_003_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (11),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (pll_c2_out),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_ext),                               //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src4_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src4_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src4_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src4_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src4_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (11),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_ext),                               //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (pll_c2_out),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	nios_simple_irq_mapper irq_mapper (
		.clk           (pll_c2_out),                         //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c3_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c2_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c3_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c2_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (pll_c3_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c2_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

endmodule
